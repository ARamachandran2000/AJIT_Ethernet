-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity AccessRegister is -- 
  generic (tag_length : integer); 
  port ( -- 
    rwbar : in  std_logic_vector(0 downto 0);
    bmask : in  std_logic_vector(3 downto 0);
    register_index : in  std_logic_vector(5 downto 0);
    wdata : in  std_logic_vector(31 downto 0);
    rdata : out  std_logic_vector(31 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity AccessRegister;
architecture AccessRegister_arch of AccessRegister is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 43)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal bmask_buffer :  std_logic_vector(3 downto 0);
  signal bmask_update_enable: Boolean;
  signal register_index_buffer :  std_logic_vector(5 downto 0);
  signal register_index_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(31 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(31 downto 0);
  signal rdata_update_enable: Boolean;
  signal AccessRegister_CP_0_start: Boolean;
  signal AccessRegister_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_req_0 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_ack_0 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_req_1 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_ack_1 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_req_0 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_ack_0 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_req_1 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "AccessRegister_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 43) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(4 downto 1) <= bmask;
  bmask_buffer <= in_buffer_data_out(4 downto 1);
  in_buffer_data_in(10 downto 5) <= register_index;
  register_index_buffer <= in_buffer_data_out(10 downto 5);
  in_buffer_data_in(42 downto 11) <= wdata;
  wdata_buffer <= in_buffer_data_out(42 downto 11);
  in_buffer_data_in(tag_length + 42 downto 43) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 42 downto 43);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  AccessRegister_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "AccessRegister_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= AccessRegister_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= AccessRegister_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= AccessRegister_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  AccessRegister_CP_0: Block -- control-path 
    signal AccessRegister_CP_0_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    AccessRegister_CP_0_elements(0) <= AccessRegister_CP_0_start;
    AccessRegister_CP_0_symbol <= AccessRegister_CP_0_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_sample_start_
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Sample/req
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/$entry
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_sample_start_
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Sample/rr
      -- 
    rr_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(0), ack => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_req_0); -- 
    req_13_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_13_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(0), ack => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_sample_completed_
      -- CP-element group 1: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_update_start_
      -- CP-element group 1: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Sample/ack
      -- CP-element group 1: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Update/$entry
      -- CP-element group 1: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Update/req
      -- 
    ack_14_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_ack_0, ack => AccessRegister_CP_0_elements(1)); -- 
    req_18_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_18_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(1), ack => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_update_completed_
      -- CP-element group 2: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Update/$exit
      -- CP-element group 2: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Update/ack
      -- 
    ack_19_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_ack_1, ack => AccessRegister_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_sample_completed_
      -- CP-element group 3: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_update_start_
      -- CP-element group 3: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Sample/ra
      -- CP-element group 3: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Update/$entry
      -- CP-element group 3: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Update/cr
      -- 
    ra_28_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_ack_0, ack => AccessRegister_CP_0_elements(3)); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(3), ack => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_update_completed_
      -- CP-element group 4: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Update/$exit
      -- CP-element group 4: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Update/ca
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_ack_1, ack => AccessRegister_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_77_to_assign_stmt_95/$exit
      -- 
    AccessRegister_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "AccessRegister_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= AccessRegister_CP_0_elements(4) & AccessRegister_CP_0_elements(2);
      gj_AccessRegister_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => AccessRegister_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u5_72_wire : std_logic_vector(4 downto 0);
    signal CONCAT_u6_u38_75_wire : std_logic_vector(37 downto 0);
    signal request_77 : std_logic_vector(42 downto 0);
    signal response_89 : std_logic_vector(32 downto 0);
    -- 
  begin -- 
    -- flow-through slice operator slice_94_inst
    rdata_buffer <= response_89(31 downto 0);
    -- binary operator CONCAT_u1_u5_72_inst
    process(rwbar_buffer, bmask_buffer) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApConcat_proc(rwbar_buffer, bmask_buffer, tmp_var);
      CONCAT_u1_u5_72_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u5_u43_76_inst
    process(CONCAT_u1_u5_72_wire, CONCAT_u6_u38_75_wire) -- 
      variable tmp_var : std_logic_vector(42 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u5_72_wire, CONCAT_u6_u38_75_wire, tmp_var);
      request_77 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u6_u38_75_inst
    process(register_index_buffer, wdata_buffer) -- 
      variable tmp_var : std_logic_vector(37 downto 0); -- 
    begin -- 
      ApConcat_proc(register_index_buffer, wdata_buffer, tmp_var);
      CONCAT_u6_u38_75_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_req_0;
      RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_req_1;
      RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      response_89 <= data_out(32 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0_gI: SplitGuardInterface generic map(name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0: InputPortRevised -- 
        generic map ( name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req(0),
          oack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack(0),
          odata => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_req_0;
      WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_req_1;
      WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= request_77;
      NIC_REQUEST_REGISTER_ACCESS_PIPE_write_0_gI: SplitGuardInterface generic map(name => "NIC_REQUEST_REGISTER_ACCESS_PIPE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_REQUEST_REGISTER_ACCESS_PIPE_write_0: OutputPortRevised -- 
        generic map ( name => "NIC_REQUEST_REGISTER_ACCESS_PIPE", data_width => 43, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req(0),
          oack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack(0),
          odata => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data(42 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end AccessRegister_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity NicRegisterAccessDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(42 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(32 downto 0);
    UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
    UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
    UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
    UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity NicRegisterAccessDaemon;
architecture NicRegisterAccessDaemon_arch of NicRegisterAccessDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal NicRegisterAccessDaemon_CP_116_start: Boolean;
  signal NicRegisterAccessDaemon_CP_116_symbol: Boolean;
  -- volatile/operator module components. 
  component UpdateRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      bmask : in  std_logic_vector(3 downto 0);
      rval : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      index : in  std_logic_vector(5 downto 0);
      wval : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal do_while_stmt_179_branch_req_0 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_req_0 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_ack_0 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_req_1 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_ack_1 : boolean;
  signal array_obj_ref_203_load_0_req_0 : boolean;
  signal array_obj_ref_203_load_0_ack_0 : boolean;
  signal array_obj_ref_203_load_0_req_1 : boolean;
  signal array_obj_ref_203_load_0_ack_1 : boolean;
  signal W_rwbar_212_delayed_5_0_208_inst_req_0 : boolean;
  signal W_rwbar_212_delayed_5_0_208_inst_ack_0 : boolean;
  signal W_rwbar_212_delayed_5_0_208_inst_req_1 : boolean;
  signal W_rwbar_212_delayed_5_0_208_inst_ack_1 : boolean;
  signal W_bmask_213_delayed_5_0_211_inst_req_0 : boolean;
  signal W_bmask_213_delayed_5_0_211_inst_ack_0 : boolean;
  signal W_bmask_213_delayed_5_0_211_inst_req_1 : boolean;
  signal W_bmask_213_delayed_5_0_211_inst_ack_1 : boolean;
  signal W_wdata_215_delayed_5_0_214_inst_req_0 : boolean;
  signal W_wdata_215_delayed_5_0_214_inst_ack_0 : boolean;
  signal W_wdata_215_delayed_5_0_214_inst_req_1 : boolean;
  signal W_wdata_215_delayed_5_0_214_inst_ack_1 : boolean;
  signal W_index_216_delayed_5_0_217_inst_req_0 : boolean;
  signal W_index_216_delayed_5_0_217_inst_ack_0 : boolean;
  signal W_index_216_delayed_5_0_217_inst_req_1 : boolean;
  signal W_index_216_delayed_5_0_217_inst_ack_1 : boolean;
  signal call_stmt_226_call_req_0 : boolean;
  signal call_stmt_226_call_ack_0 : boolean;
  signal call_stmt_226_call_req_1 : boolean;
  signal call_stmt_226_call_ack_1 : boolean;
  signal W_rwbar_220_delayed_5_0_227_inst_req_0 : boolean;
  signal W_rwbar_220_delayed_5_0_227_inst_ack_0 : boolean;
  signal W_rwbar_220_delayed_5_0_227_inst_req_1 : boolean;
  signal W_rwbar_220_delayed_5_0_227_inst_ack_1 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_req_0 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_ack_0 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_req_1 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_ack_1 : boolean;
  signal do_while_stmt_179_branch_ack_0 : boolean;
  signal do_while_stmt_179_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "NicRegisterAccessDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  NicRegisterAccessDaemon_CP_116_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "NicRegisterAccessDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= NicRegisterAccessDaemon_CP_116_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= NicRegisterAccessDaemon_CP_116_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= NicRegisterAccessDaemon_CP_116_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  NicRegisterAccessDaemon_CP_116: Block -- control-path 
    signal NicRegisterAccessDaemon_CP_116_elements: BooleanArray(50 downto 0);
    -- 
  begin -- 
    NicRegisterAccessDaemon_CP_116_elements(0) <= NicRegisterAccessDaemon_CP_116_start;
    NicRegisterAccessDaemon_CP_116_symbol <= NicRegisterAccessDaemon_CP_116_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_178/$entry
      -- CP-element group 0: 	 branch_block_stmt_178/branch_block_stmt_178__entry__
      -- CP-element group 0: 	 branch_block_stmt_178/do_while_stmt_179__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	50 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_178/$exit
      -- CP-element group 1: 	 branch_block_stmt_178/branch_block_stmt_178__exit__
      -- CP-element group 1: 	 branch_block_stmt_178/do_while_stmt_179__exit__
      -- 
    NicRegisterAccessDaemon_CP_116_elements(1) <= NicRegisterAccessDaemon_CP_116_elements(50);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_178/do_while_stmt_179/$entry
      -- CP-element group 2: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179__entry__
      -- 
    NicRegisterAccessDaemon_CP_116_elements(2) <= NicRegisterAccessDaemon_CP_116_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	50 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179__exit__
      -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_178/do_while_stmt_179/loop_back
      -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	45 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	48 
    -- CP-element group 5: 	49 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_178/do_while_stmt_179/condition_done
      -- CP-element group 5: 	 branch_block_stmt_178/do_while_stmt_179/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_178/do_while_stmt_179/loop_taken/$entry
      -- 
    NicRegisterAccessDaemon_CP_116_elements(5) <= NicRegisterAccessDaemon_CP_116_elements(45);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	47 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_178/do_while_stmt_179/loop_body_done
      -- 
    NicRegisterAccessDaemon_CP_116_elements(6) <= NicRegisterAccessDaemon_CP_116_elements(47);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/back_edge_to_loop_body
      -- 
    NicRegisterAccessDaemon_CP_116_elements(7) <= NicRegisterAccessDaemon_CP_116_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/first_time_through_loop_body
      -- 
    NicRegisterAccessDaemon_CP_116_elements(8) <= NicRegisterAccessDaemon_CP_116_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	45 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/loop_body_start
      -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	13 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Sample/rr
      -- 
    rr_149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(10), ack => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(9) & NicRegisterAccessDaemon_CP_116_elements(13);
      gj_NicRegisterAccessDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	20 
    -- CP-element group 11: 	24 
    -- CP-element group 11: 	28 
    -- CP-element group 11: 	32 
    -- CP-element group 11: 	40 
    -- CP-element group 11: 	16 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_update_start_
      -- CP-element group 11: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Update/cr
      -- 
    cr_154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(11), ack => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(12) & NicRegisterAccessDaemon_CP_116_elements(20) & NicRegisterAccessDaemon_CP_116_elements(24) & NicRegisterAccessDaemon_CP_116_elements(28) & NicRegisterAccessDaemon_CP_116_elements(32) & NicRegisterAccessDaemon_CP_116_elements(40) & NicRegisterAccessDaemon_CP_116_elements(16);
      gj_NicRegisterAccessDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Sample/ra
      -- 
    ra_150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	18 
    -- CP-element group 13: 	22 
    -- CP-element group 13: 	26 
    -- CP-element group 13: 	30 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	14 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	10 
    -- CP-element group 13:  members (29) 
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_resize_0/$entry
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_resize_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_resize_0/index_resize_req
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_resize_0/index_resize_ack
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_scale_0/$entry
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_scale_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_scale_0/scale_rename_req
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_scale_0/scale_rename_ack
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_final_index_sum_regn/$entry
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_final_index_sum_regn/$exit
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_final_index_sum_regn/req
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_final_index_sum_regn/ack
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_word_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_root_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_offset_calculated
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_resized_0
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_scaled_0
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_computed_0
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_base_plus_offset/$entry
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_base_plus_offset/$exit
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_base_plus_offset/sum_rename_req
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_base_plus_offset/sum_rename_ack
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_word_addrgen/$entry
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_word_addrgen/$exit
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_word_addrgen/root_register_req
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_word_addrgen/root_register_ack
      -- 
    ca_155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/word_access_start/$entry
      -- CP-element group 14: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/word_access_start/word_0/$entry
      -- CP-element group 14: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/word_access_start/word_0/rr
      -- 
    rr_201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(14), ack => array_obj_ref_203_load_0_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(37) & NicRegisterAccessDaemon_CP_116_elements(16);
      gj_NicRegisterAccessDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	36 
    -- CP-element group 15: 	43 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_update_start_
      -- CP-element group 15: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/word_access_complete/$entry
      -- CP-element group 15: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/word_access_complete/word_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/word_access_complete/word_0/cr
      -- 
    cr_212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(15), ack => array_obj_ref_203_load_0_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(36) & NicRegisterAccessDaemon_CP_116_elements(43);
      gj_NicRegisterAccessDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	46 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/word_access_start/$exit
      -- CP-element group 16: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/word_access_start/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/word_access_start/word_0/ra
      -- 
    ra_202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_203_load_0_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	34 
    -- CP-element group 17: 	42 
    -- CP-element group 17:  members (9) 
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/word_access_complete/$exit
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/word_access_complete/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/word_access_complete/word_0/ca
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/array_obj_ref_203_Merge/$entry
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/array_obj_ref_203_Merge/$exit
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/array_obj_ref_203_Merge/merge_req
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/array_obj_ref_203_Merge/merge_ack
      -- 
    ca_213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_203_load_0_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	13 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Sample/req
      -- 
    req_226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(18), ack => W_rwbar_212_delayed_5_0_208_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(20);
      gj_NicRegisterAccessDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	36 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_update_start_
      -- CP-element group 19: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Update/req
      -- 
    req_231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(19), ack => W_rwbar_212_delayed_5_0_208_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(36);
      gj_NicRegisterAccessDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: 	11 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Sample/ack
      -- 
    ack_227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_212_delayed_5_0_208_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	34 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Update/ack
      -- 
    ack_232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_212_delayed_5_0_208_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	13 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Sample/req
      -- 
    req_240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(22), ack => W_bmask_213_delayed_5_0_211_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(24);
      gj_NicRegisterAccessDaemon_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	36 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_update_start_
      -- CP-element group 23: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Update/req
      -- 
    req_245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(23), ack => W_bmask_213_delayed_5_0_211_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(36);
      gj_NicRegisterAccessDaemon_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: 	11 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Sample/ack
      -- 
    ack_241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_213_delayed_5_0_211_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	34 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Update/ack
      -- 
    ack_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_213_delayed_5_0_211_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(25)); -- 
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	13 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Sample/req
      -- 
    req_254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(26), ack => W_wdata_215_delayed_5_0_214_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(28);
      gj_NicRegisterAccessDaemon_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	36 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_update_start_
      -- CP-element group 27: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Update/req
      -- 
    req_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(27), ack => W_wdata_215_delayed_5_0_214_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(36);
      gj_NicRegisterAccessDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: 	11 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Sample/ack
      -- 
    ack_255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_215_delayed_5_0_214_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	34 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Update/ack
      -- 
    ack_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_215_delayed_5_0_214_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(29)); -- 
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	13 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Sample/req
      -- 
    req_268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(30), ack => W_index_216_delayed_5_0_217_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(32);
      gj_NicRegisterAccessDaemon_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	36 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_update_start_
      -- CP-element group 31: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Update/req
      -- 
    req_273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(31), ack => W_index_216_delayed_5_0_217_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(36);
      gj_NicRegisterAccessDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: 	11 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Sample/ack
      -- 
    ack_269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_216_delayed_5_0_217_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Update/ack
      -- 
    ack_274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_216_delayed_5_0_217_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(33)); -- 
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	17 
    -- CP-element group 34: 	21 
    -- CP-element group 34: 	25 
    -- CP-element group 34: 	29 
    -- CP-element group 34: 	33 
    -- CP-element group 34: 	46 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Sample/crr
      -- 
    crr_282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(34), ack => call_stmt_226_call_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 31,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(17) & NicRegisterAccessDaemon_CP_116_elements(21) & NicRegisterAccessDaemon_CP_116_elements(25) & NicRegisterAccessDaemon_CP_116_elements(29) & NicRegisterAccessDaemon_CP_116_elements(33) & NicRegisterAccessDaemon_CP_116_elements(46) & NicRegisterAccessDaemon_CP_116_elements(36);
      gj_NicRegisterAccessDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_update_start_
      -- CP-element group 35: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Update/ccr
      -- 
    ccr_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(35), ack => call_stmt_226_call_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(37);
      gj_NicRegisterAccessDaemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	19 
    -- CP-element group 36: 	23 
    -- CP-element group 36: 	27 
    -- CP-element group 36: 	31 
    -- CP-element group 36: 	34 
    -- CP-element group 36: 	15 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Sample/cra
      -- 
    cra_283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_226_call_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(36)); -- 
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	47 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: 	14 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Update/cca
      -- CP-element group 37: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/ring_reenable_memory_space_0
      -- 
    cca_288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_226_call_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	40 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Sample/req
      -- 
    req_296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(38), ack => W_rwbar_220_delayed_5_0_227_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(40);
      gj_NicRegisterAccessDaemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	43 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_update_start_
      -- CP-element group 39: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Update/req
      -- 
    req_301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(39), ack => W_rwbar_220_delayed_5_0_227_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(43);
      gj_NicRegisterAccessDaemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: 	11 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Sample/ack
      -- 
    ack_297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_220_delayed_5_0_227_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Update/ack
      -- 
    ack_302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_220_delayed_5_0_227_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	17 
    -- CP-element group 42: 	41 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Sample/req
      -- 
    req_310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(42), ack => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(17) & NicRegisterAccessDaemon_CP_116_elements(41) & NicRegisterAccessDaemon_CP_116_elements(44);
      gj_NicRegisterAccessDaemon_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	39 
    -- CP-element group 43: 	15 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_update_start_
      -- CP-element group 43: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Update/req
      -- 
    ack_311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(43)); -- 
    req_315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(43), ack => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_req_1); -- 
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	47 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Update/ack
      -- 
    ack_316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(44)); -- 
    -- CP-element group 45:  transition  output  delay-element  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	9 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	5 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/condition_evaluated
      -- CP-element group 45: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/loop_body_delay_to_condition_start
      -- 
    condition_evaluated_140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(45), ack => do_while_stmt_179_branch_req_0); -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(45) is a control-delay.
    cp_element_45_delay: control_delay_element  generic map(name => " 45_delay", delay_value => 1)  port map(req => NicRegisterAccessDaemon_CP_116_elements(9), ack => NicRegisterAccessDaemon_CP_116_elements(45), clk => clk, reset =>reset);
    -- CP-element group 46:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	16 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	34 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_call_stmt_226_delay
      -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(46) is a control-delay.
    cp_element_46_delay: control_delay_element  generic map(name => " 46_delay", delay_value => 1)  port map(req => NicRegisterAccessDaemon_CP_116_elements(16), ack => NicRegisterAccessDaemon_CP_116_elements(46), clk => clk, reset =>reset);
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	37 
    -- CP-element group 47: 	44 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	6 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/$exit
      -- 
    NicRegisterAccessDaemon_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(37) & NicRegisterAccessDaemon_CP_116_elements(44);
      gj_NicRegisterAccessDaemon_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	5 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_178/do_while_stmt_179/loop_exit/$exit
      -- CP-element group 48: 	 branch_block_stmt_178/do_while_stmt_179/loop_exit/ack
      -- 
    ack_323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_179_branch_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	5 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_178/do_while_stmt_179/loop_taken/$exit
      -- CP-element group 49: 	 branch_block_stmt_178/do_while_stmt_179/loop_taken/ack
      -- 
    ack_327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_179_branch_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(49)); -- 
    -- CP-element group 50:  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	3 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	1 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_178/do_while_stmt_179/$exit
      -- 
    NicRegisterAccessDaemon_CP_116_elements(50) <= NicRegisterAccessDaemon_CP_116_elements(3);
    NicRegisterAccessDaemon_do_while_stmt_179_terminator_328: loop_terminator -- 
      generic map (name => " NicRegisterAccessDaemon_do_while_stmt_179_terminator_328", max_iterations_in_flight =>31) 
      port map(loop_body_exit => NicRegisterAccessDaemon_CP_116_elements(6),loop_continue => NicRegisterAccessDaemon_CP_116_elements(49),loop_terminate => NicRegisterAccessDaemon_CP_116_elements(48),loop_back => NicRegisterAccessDaemon_CP_116_elements(4),loop_exit => NicRegisterAccessDaemon_CP_116_elements(3),clk => clk, reset => reset); -- 
    entry_tmerge_141_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= NicRegisterAccessDaemon_CP_116_elements(7);
        preds(1)  <= NicRegisterAccessDaemon_CP_116_elements(8);
        entry_tmerge_141 : transition_merge -- 
          generic map(name => " entry_tmerge_141")
          port map (preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_index_202_resized : std_logic_vector(5 downto 0);
    signal R_index_202_scaled : std_logic_vector(5 downto 0);
    signal array_obj_ref_203_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_203_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_203_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_203_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_203_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_203_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_203_word_offset_0 : std_logic_vector(5 downto 0);
    signal bmask_192 : std_logic_vector(3 downto 0);
    signal bmask_213_delayed_5_0_213 : std_logic_vector(3 downto 0);
    signal index_196 : std_logic_vector(5 downto 0);
    signal index_216_delayed_5_0_219 : std_logic_vector(5 downto 0);
    signal konst_247_wire_constant : std_logic_vector(0 downto 0);
    signal rdata_236 : std_logic_vector(31 downto 0);
    signal req_183 : std_logic_vector(42 downto 0);
    signal resp_242 : std_logic_vector(32 downto 0);
    signal rval_204 : std_logic_vector(31 downto 0);
    signal rwbar_188 : std_logic_vector(0 downto 0);
    signal rwbar_212_delayed_5_0_210 : std_logic_vector(0 downto 0);
    signal rwbar_220_delayed_5_0_229 : std_logic_vector(0 downto 0);
    signal type_cast_234_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_239_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_200 : std_logic_vector(31 downto 0);
    signal wdata_215_delayed_5_0_216 : std_logic_vector(31 downto 0);
    signal wval_226 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_203_offset_scale_factor_0 <= "000001";
    array_obj_ref_203_resized_base_address <= "000000";
    array_obj_ref_203_word_offset_0 <= "000000";
    konst_247_wire_constant <= "1";
    type_cast_234_wire_constant <= "00000000000000000000000000000000";
    type_cast_239_wire_constant <= "0";
    -- flow-through select operator MUX_235_inst
    rdata_236 <= rval_204 when (rwbar_220_delayed_5_0_229(0) /=  '0') else type_cast_234_wire_constant;
    -- flow-through slice operator slice_187_inst
    rwbar_188 <= req_183(42 downto 42);
    -- flow-through slice operator slice_191_inst
    bmask_192 <= req_183(41 downto 38);
    -- flow-through slice operator slice_195_inst
    index_196 <= req_183(37 downto 32);
    -- flow-through slice operator slice_199_inst
    wdata_200 <= req_183(31 downto 0);
    W_bmask_213_delayed_5_0_211_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_bmask_213_delayed_5_0_211_inst_req_0;
      W_bmask_213_delayed_5_0_211_inst_ack_0<= wack(0);
      rreq(0) <= W_bmask_213_delayed_5_0_211_inst_req_1;
      W_bmask_213_delayed_5_0_211_inst_ack_1<= rack(0);
      W_bmask_213_delayed_5_0_211_inst : InterlockBuffer generic map ( -- 
        name => "W_bmask_213_delayed_5_0_211_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => bmask_192,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => bmask_213_delayed_5_0_213,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_index_216_delayed_5_0_217_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_index_216_delayed_5_0_217_inst_req_0;
      W_index_216_delayed_5_0_217_inst_ack_0<= wack(0);
      rreq(0) <= W_index_216_delayed_5_0_217_inst_req_1;
      W_index_216_delayed_5_0_217_inst_ack_1<= rack(0);
      W_index_216_delayed_5_0_217_inst : InterlockBuffer generic map ( -- 
        name => "W_index_216_delayed_5_0_217_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => index_196,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => index_216_delayed_5_0_219,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_212_delayed_5_0_208_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_212_delayed_5_0_208_inst_req_0;
      W_rwbar_212_delayed_5_0_208_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_212_delayed_5_0_208_inst_req_1;
      W_rwbar_212_delayed_5_0_208_inst_ack_1<= rack(0);
      W_rwbar_212_delayed_5_0_208_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_212_delayed_5_0_208_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_212_delayed_5_0_210,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_220_delayed_5_0_227_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_220_delayed_5_0_227_inst_req_0;
      W_rwbar_220_delayed_5_0_227_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_220_delayed_5_0_227_inst_req_1;
      W_rwbar_220_delayed_5_0_227_inst_ack_1<= rack(0);
      W_rwbar_220_delayed_5_0_227_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_220_delayed_5_0_227_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_220_delayed_5_0_229,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_wdata_215_delayed_5_0_214_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_wdata_215_delayed_5_0_214_inst_req_0;
      W_wdata_215_delayed_5_0_214_inst_ack_0<= wack(0);
      rreq(0) <= W_wdata_215_delayed_5_0_214_inst_req_1;
      W_wdata_215_delayed_5_0_214_inst_ack_1<= rack(0);
      W_wdata_215_delayed_5_0_214_inst : InterlockBuffer generic map ( -- 
        name => "W_wdata_215_delayed_5_0_214_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => wdata_200,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => wdata_215_delayed_5_0_216,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_203_addr_0
    process(array_obj_ref_203_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_203_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_203_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_203_gather_scatter
    process(array_obj_ref_203_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_203_data_0;
      ov(31 downto 0) := iv;
      rval_204 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_203_index_0_rename
    process(R_index_202_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_202_resized;
      ov(5 downto 0) := iv;
      R_index_202_scaled <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_203_index_0_resize
    process(index_196) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_196;
      ov(5 downto 0) := iv;
      R_index_202_resized <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_203_index_offset
    process(R_index_202_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_202_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_203_final_offset <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_203_root_address_inst
    process(array_obj_ref_203_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_203_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_203_root_address <= ov(5 downto 0);
      --
    end process;
    do_while_stmt_179_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_247_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_179_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_179_branch_req_0,
          ack0 => do_while_stmt_179_branch_ack_0,
          ack1 => do_while_stmt_179_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u1_u33_241_inst
    process(type_cast_239_wire_constant, rdata_236) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_239_wire_constant, rdata_236, tmp_var);
      resp_242 <= tmp_var; --
    end process;
    -- shared load operator group (0) : array_obj_ref_203_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_203_load_0_req_0;
      array_obj_ref_203_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_203_load_0_req_1;
      array_obj_ref_203_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_203_word_address_0;
      array_obj_ref_203_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 6,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(5 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(42 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_req_0;
      RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_req_1;
      RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      req_183 <= data_out(42 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0_gI: SplitGuardInterface generic map(name => "NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0: InputPortRevised -- 
        generic map ( name => "NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0", data_width => 43,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req(0),
          oack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack(0),
          odata => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data(42 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_req_0;
      WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_req_1;
      WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= resp_242;
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_write_0_gI: SplitGuardInterface generic map(name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_write_0: OutputPortRevised -- 
        generic map ( name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req(0),
          oack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack(0),
          odata => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_226_call 
    UpdateRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(73 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_226_call_req_0;
      call_stmt_226_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_226_call_req_1;
      call_stmt_226_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not rwbar_212_delayed_5_0_210(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      UpdateRegister_call_group_0_gI: SplitGuardInterface generic map(name => "UpdateRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= bmask_213_delayed_5_0_213 & rval_204 & wdata_215_delayed_5_0_216 & index_216_delayed_5_0_219;
      wval_226 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 74,
        owidth => 74,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => UpdateRegister_call_reqs(0),
          ackR => UpdateRegister_call_acks(0),
          dataR => UpdateRegister_call_data(73 downto 0),
          tagR => UpdateRegister_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => UpdateRegister_return_acks(0), -- cross-over
          ackL => UpdateRegister_return_reqs(0), -- cross-over
          dataL => UpdateRegister_return_data(31 downto 0),
          tagL => UpdateRegister_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end NicRegisterAccessDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity ReceiveEngineDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    FREE_Q : in std_logic_vector(35 downto 0);
    CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
    populateRxQueue_call_reqs : out  std_logic_vector(0 downto 0);
    populateRxQueue_call_acks : in   std_logic_vector(0 downto 0);
    populateRxQueue_call_data : out  std_logic_vector(35 downto 0);
    populateRxQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    populateRxQueue_return_reqs : out  std_logic_vector(0 downto 0);
    populateRxQueue_return_acks : in   std_logic_vector(0 downto 0);
    populateRxQueue_return_tag :  in   std_logic_vector(0 downto 0);
    popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_call_data : out  std_logic_vector(36 downto 0);
    popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_return_data : in   std_logic_vector(32 downto 0);
    popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
    loadBuffer_call_reqs : out  std_logic_vector(0 downto 0);
    loadBuffer_call_acks : in   std_logic_vector(0 downto 0);
    loadBuffer_call_data : out  std_logic_vector(35 downto 0);
    loadBuffer_call_tag  :  out  std_logic_vector(0 downto 0);
    loadBuffer_return_reqs : out  std_logic_vector(0 downto 0);
    loadBuffer_return_acks : in   std_logic_vector(0 downto 0);
    loadBuffer_return_data : in   std_logic_vector(0 downto 0);
    loadBuffer_return_tag :  in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity ReceiveEngineDaemon;
architecture ReceiveEngineDaemon_arch of ReceiveEngineDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ReceiveEngineDaemon_CP_1640_start: Boolean;
  signal ReceiveEngineDaemon_CP_1640_symbol: Boolean;
  -- volatile/operator module components. 
  component populateRxQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
      NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(67 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(31 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadBuffer is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_data : out  std_logic_vector(51 downto 0);
      writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_data : out  std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_data : in   std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_data : out  std_logic_vector(71 downto 0);
      writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_return_data : in   std_logic_vector(16 downto 0);
      writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_inst_req_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_inst_ack_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_inst_req_1 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_inst_ack_1 : boolean;
  signal if_stmt_971_branch_req_0 : boolean;
  signal if_stmt_971_branch_ack_1 : boolean;
  signal if_stmt_971_branch_ack_0 : boolean;
  signal do_while_stmt_979_branch_req_0 : boolean;
  signal call_stmt_987_call_req_0 : boolean;
  signal call_stmt_987_call_ack_0 : boolean;
  signal call_stmt_987_call_req_1 : boolean;
  signal call_stmt_987_call_ack_1 : boolean;
  signal call_stmt_1005_call_req_0 : boolean;
  signal call_stmt_1005_call_ack_0 : boolean;
  signal call_stmt_1005_call_req_1 : boolean;
  signal call_stmt_1005_call_ack_1 : boolean;
  signal NOT_u1_u1_1008_inst_req_0 : boolean;
  signal NOT_u1_u1_1008_inst_ack_0 : boolean;
  signal NOT_u1_u1_1008_inst_req_1 : boolean;
  signal NOT_u1_u1_1008_inst_ack_1 : boolean;
  signal NOT_u1_u1_1018_inst_req_0 : boolean;
  signal NOT_u1_u1_1018_inst_ack_0 : boolean;
  signal NOT_u1_u1_1018_inst_req_1 : boolean;
  signal NOT_u1_u1_1018_inst_ack_1 : boolean;
  signal W_rx_buffer_pointer_36_1016_delayed_10_0_1034_inst_req_0 : boolean;
  signal W_rx_buffer_pointer_36_1016_delayed_10_0_1034_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_36_1016_delayed_10_0_1034_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_36_1016_delayed_10_0_1034_inst_ack_1 : boolean;
  signal call_stmt_1039_call_req_0 : boolean;
  signal call_stmt_1039_call_ack_0 : boolean;
  signal call_stmt_1039_call_req_1 : boolean;
  signal call_stmt_1039_call_ack_1 : boolean;
  signal W_rx_buffer_pointer_36_1024_delayed_10_0_1042_inst_req_0 : boolean;
  signal W_rx_buffer_pointer_36_1024_delayed_10_0_1042_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_36_1024_delayed_10_0_1042_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_36_1024_delayed_10_0_1042_inst_ack_1 : boolean;
  signal call_stmt_1052_call_req_0 : boolean;
  signal call_stmt_1052_call_ack_0 : boolean;
  signal call_stmt_1052_call_req_1 : boolean;
  signal call_stmt_1052_call_ack_1 : boolean;
  signal do_while_stmt_979_branch_ack_0 : boolean;
  signal do_while_stmt_979_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "ReceiveEngineDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  ReceiveEngineDaemon_CP_1640_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "ReceiveEngineDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_1640_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_1640_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_1640_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  ReceiveEngineDaemon_CP_1640: Block -- control-path 
    signal ReceiveEngineDaemon_CP_1640_elements: BooleanArray(51 downto 0);
    -- 
  begin -- 
    ReceiveEngineDaemon_CP_1640_elements(0) <= ReceiveEngineDaemon_CP_1640_start;
    ReceiveEngineDaemon_CP_1640_symbol <= ReceiveEngineDaemon_CP_1640_elements(3);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_967/$entry
      -- CP-element group 0: 	 assign_stmt_967/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_sample_start_
      -- CP-element group 0: 	 assign_stmt_967/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_967/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_Sample/req
      -- 
    req_1653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(0), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_967/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_sample_completed_
      -- CP-element group 1: 	 assign_stmt_967/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_update_start_
      -- CP-element group 1: 	 assign_stmt_967/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_967/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_Sample/ack
      -- CP-element group 1: 	 assign_stmt_967/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_Update/$entry
      -- CP-element group 1: 	 assign_stmt_967/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_Update/req
      -- 
    ack_1654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_inst_ack_0, ack => ReceiveEngineDaemon_CP_1640_elements(1)); -- 
    req_1658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(1), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_inst_req_1); -- 
    -- CP-element group 2:  branch  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	51 
    -- CP-element group 2:  members (10) 
      -- CP-element group 2: 	 assign_stmt_967/$exit
      -- CP-element group 2: 	 assign_stmt_967/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_update_completed_
      -- CP-element group 2: 	 assign_stmt_967/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_Update/$exit
      -- CP-element group 2: 	 assign_stmt_967/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_Update/ack
      -- CP-element group 2: 	 branch_block_stmt_968/$entry
      -- CP-element group 2: 	 branch_block_stmt_968/branch_block_stmt_968__entry__
      -- CP-element group 2: 	 branch_block_stmt_968/merge_stmt_970__entry__
      -- CP-element group 2: 	 branch_block_stmt_968/merge_stmt_970_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_968/merge_stmt_970__entry___PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_968/merge_stmt_970__entry___PhiReq/$exit
      -- 
    ack_1659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_inst_ack_1, ack => ReceiveEngineDaemon_CP_1640_elements(2)); -- 
    -- CP-element group 3:  transition  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 $exit
      -- CP-element group 3: 	 branch_block_stmt_968/$exit
      -- CP-element group 3: 	 branch_block_stmt_968/branch_block_stmt_968__exit__
      -- 
    ReceiveEngineDaemon_CP_1640_elements(3) <= false; 
    -- CP-element group 4:  transition  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	50 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	51 
    -- CP-element group 4:  members (4) 
      -- CP-element group 4: 	 branch_block_stmt_968/do_while_stmt_979__exit__
      -- CP-element group 4: 	 branch_block_stmt_968/disable_loopback
      -- CP-element group 4: 	 branch_block_stmt_968/disable_loopback_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_968/disable_loopback_PhiReq/$exit
      -- 
    ReceiveEngineDaemon_CP_1640_elements(4) <= ReceiveEngineDaemon_CP_1640_elements(50);
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	51 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	51 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_968/if_stmt_971_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_968/if_stmt_971_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_968/not_enabled_yet_loopback
      -- CP-element group 5: 	 branch_block_stmt_968/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_968/not_enabled_yet_loopback_PhiReq/$exit
      -- 
    if_choice_transition_1732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_971_branch_ack_1, ack => ReceiveEngineDaemon_CP_1640_elements(5)); -- 
    -- CP-element group 6:  merge  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	51 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (4) 
      -- CP-element group 6: 	 branch_block_stmt_968/if_stmt_971__exit__
      -- CP-element group 6: 	 branch_block_stmt_968/do_while_stmt_979__entry__
      -- CP-element group 6: 	 branch_block_stmt_968/if_stmt_971_else_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_968/if_stmt_971_else_link/else_choice_transition
      -- 
    else_choice_transition_1736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_971_branch_ack_0, ack => ReceiveEngineDaemon_CP_1640_elements(6)); -- 
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_968/do_while_stmt_979/$entry
      -- CP-element group 7: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979__entry__
      -- 
    ReceiveEngineDaemon_CP_1640_elements(7) <= ReceiveEngineDaemon_CP_1640_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	50 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979__exit__
      -- 
    -- Element group ReceiveEngineDaemon_CP_1640_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_968/do_while_stmt_979/loop_back
      -- 
    -- Element group ReceiveEngineDaemon_CP_1640_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	47 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	48 
    -- CP-element group 10: 	49 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_968/do_while_stmt_979/condition_done
      -- CP-element group 10: 	 branch_block_stmt_968/do_while_stmt_979/loop_exit/$entry
      -- CP-element group 10: 	 branch_block_stmt_968/do_while_stmt_979/loop_taken/$entry
      -- 
    ReceiveEngineDaemon_CP_1640_elements(10) <= ReceiveEngineDaemon_CP_1640_elements(47);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	46 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_968/do_while_stmt_979/loop_body_done
      -- 
    ReceiveEngineDaemon_CP_1640_elements(11) <= ReceiveEngineDaemon_CP_1640_elements(46);
    -- CP-element group 12:  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/back_edge_to_loop_body
      -- 
    ReceiveEngineDaemon_CP_1640_elements(12) <= ReceiveEngineDaemon_CP_1640_elements(9);
    -- CP-element group 13:  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/first_time_through_loop_body
      -- 
    ReceiveEngineDaemon_CP_1640_elements(13) <= ReceiveEngineDaemon_CP_1640_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	47 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/$entry
      -- CP-element group 14: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/loop_body_start
      -- 
    -- Element group ReceiveEngineDaemon_CP_1640_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	46 
    -- CP-element group 15: 	17 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_987_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_987_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_987_Sample/crr
      -- 
    crr_1761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(15), ack => call_stmt_987_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1640_elements(14) & ReceiveEngineDaemon_CP_1640_elements(46) & ReceiveEngineDaemon_CP_1640_elements(17);
      gj_ReceiveEngineDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1640_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	41 
    -- CP-element group 16: 	46 
    -- CP-element group 16: 	25 
    -- CP-element group 16: 	21 
    -- CP-element group 16: 	29 
    -- CP-element group 16: 	33 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_987_update_start_
      -- CP-element group 16: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_987_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_987_Update/ccr
      -- 
    ccr_1766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(16), ack => call_stmt_987_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1640_elements(41) & ReceiveEngineDaemon_CP_1640_elements(46) & ReceiveEngineDaemon_CP_1640_elements(25) & ReceiveEngineDaemon_CP_1640_elements(21) & ReceiveEngineDaemon_CP_1640_elements(29) & ReceiveEngineDaemon_CP_1640_elements(33);
      gj_ReceiveEngineDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1640_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	15 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_987_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_987_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_987_Sample/cra
      -- 
    cra_1762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_987_call_ack_0, ack => ReceiveEngineDaemon_CP_1640_elements(17)); -- 
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	39 
    -- CP-element group 18: 	31 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	27 
    -- CP-element group 18: 	23 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_987_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_987_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_987_Update/cca
      -- 
    cca_1767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_987_call_ack_1, ack => ReceiveEngineDaemon_CP_1640_elements(18)); -- 
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	21 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1005_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1005_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1005_Sample/crr
      -- 
    crr_1775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(19), ack => call_stmt_1005_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1640_elements(18) & ReceiveEngineDaemon_CP_1640_elements(21);
      gj_ReceiveEngineDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1640_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	37 
    -- CP-element group 20: 	45 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1005_update_start_
      -- CP-element group 20: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1005_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1005_Update/ccr
      -- 
    ccr_1780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(20), ack => call_stmt_1005_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1640_elements(37) & ReceiveEngineDaemon_CP_1640_elements(45);
      gj_ReceiveEngineDaemon_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1640_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: 	19 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1005_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1005_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1005_Sample/cra
      -- 
    cra_1776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1005_call_ack_0, ack => ReceiveEngineDaemon_CP_1640_elements(21)); -- 
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	35 
    -- CP-element group 22: 	43 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1005_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1005_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1005_Update/cca
      -- 
    cca_1781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1005_call_ack_1, ack => ReceiveEngineDaemon_CP_1640_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	18 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1008_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1008_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1008_Sample/rr
      -- 
    rr_1789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(23), ack => NOT_u1_u1_1008_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1640_elements(18) & ReceiveEngineDaemon_CP_1640_elements(25);
      gj_ReceiveEngineDaemon_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1640_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	37 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1008_update_start_
      -- CP-element group 24: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1008_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1008_Update/cr
      -- 
    cr_1794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(24), ack => NOT_u1_u1_1008_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1640_elements(37);
      gj_ReceiveEngineDaemon_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1640_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	16 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1008_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1008_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1008_Sample/ra
      -- 
    ra_1790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1008_inst_ack_0, ack => ReceiveEngineDaemon_CP_1640_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	35 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1008_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1008_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1008_Update/ca
      -- 
    ca_1795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1008_inst_ack_1, ack => ReceiveEngineDaemon_CP_1640_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	18 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1018_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1018_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1018_Sample/rr
      -- 
    rr_1803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(27), ack => NOT_u1_u1_1018_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1640_elements(18) & ReceiveEngineDaemon_CP_1640_elements(29);
      gj_ReceiveEngineDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1640_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	45 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1018_update_start_
      -- CP-element group 28: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1018_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1018_Update/cr
      -- 
    cr_1808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(28), ack => NOT_u1_u1_1018_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1640_elements(45);
      gj_ReceiveEngineDaemon_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1640_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	16 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1018_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1018_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1018_Sample/ra
      -- 
    ra_1804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1018_inst_ack_0, ack => ReceiveEngineDaemon_CP_1640_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	43 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1018_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1018_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/NOT_u1_u1_1018_Update/ca
      -- 
    ca_1809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1018_inst_ack_1, ack => ReceiveEngineDaemon_CP_1640_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	18 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1036_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1036_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1036_Sample/req
      -- 
    req_1817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(31), ack => W_rx_buffer_pointer_36_1016_delayed_10_0_1034_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1640_elements(18) & ReceiveEngineDaemon_CP_1640_elements(33);
      gj_ReceiveEngineDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1640_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	37 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1036_update_start_
      -- CP-element group 32: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1036_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1036_Update/req
      -- 
    req_1822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(32), ack => W_rx_buffer_pointer_36_1016_delayed_10_0_1034_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1640_elements(37);
      gj_ReceiveEngineDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1640_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	16 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1036_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1036_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1036_Sample/ack
      -- 
    ack_1818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1016_delayed_10_0_1034_inst_ack_0, ack => ReceiveEngineDaemon_CP_1640_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1036_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1036_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1036_Update/ack
      -- 
    ack_1823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1016_delayed_10_0_1034_inst_ack_1, ack => ReceiveEngineDaemon_CP_1640_elements(34)); -- 
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	22 
    -- CP-element group 35: 	34 
    -- CP-element group 35: 	26 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1039_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1039_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1039_Sample/crr
      -- 
    crr_1831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(35), ack => call_stmt_1039_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1640_elements(22) & ReceiveEngineDaemon_CP_1640_elements(34) & ReceiveEngineDaemon_CP_1640_elements(26) & ReceiveEngineDaemon_CP_1640_elements(37);
      gj_ReceiveEngineDaemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1640_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	38 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1039_update_start_
      -- CP-element group 36: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1039_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1039_Update/ccr
      -- 
    ccr_1836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(36), ack => call_stmt_1039_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1640_elements(38);
      gj_ReceiveEngineDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1640_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: 	20 
    -- CP-element group 37: 	24 
    -- CP-element group 37: 	32 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1039_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1039_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1039_Sample/cra
      -- 
    cra_1832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1039_call_ack_0, ack => ReceiveEngineDaemon_CP_1640_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	36 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1039_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1039_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1039_Update/cca
      -- 
    cca_1837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1039_call_ack_1, ack => ReceiveEngineDaemon_CP_1640_elements(38)); -- 
    -- CP-element group 39:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	18 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1044_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1044_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1044_Sample/req
      -- 
    req_1845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(39), ack => W_rx_buffer_pointer_36_1024_delayed_10_0_1042_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1640_elements(18) & ReceiveEngineDaemon_CP_1640_elements(41);
      gj_ReceiveEngineDaemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1640_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	45 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1044_update_start_
      -- CP-element group 40: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1044_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1044_Update/req
      -- 
    req_1850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(40), ack => W_rx_buffer_pointer_36_1024_delayed_10_0_1042_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1640_elements(45);
      gj_ReceiveEngineDaemon_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1640_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: 	16 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1044_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1044_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1044_Sample/ack
      -- 
    ack_1846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1024_delayed_10_0_1042_inst_ack_0, ack => ReceiveEngineDaemon_CP_1640_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1044_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1044_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/assign_stmt_1044_Update/ack
      -- 
    ack_1851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1024_delayed_10_0_1042_inst_ack_1, ack => ReceiveEngineDaemon_CP_1640_elements(42)); -- 
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	42 
    -- CP-element group 43: 	22 
    -- CP-element group 43: 	30 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	45 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1052_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1052_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1052_Sample/crr
      -- 
    crr_1859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(43), ack => call_stmt_1052_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1640_elements(38) & ReceiveEngineDaemon_CP_1640_elements(42) & ReceiveEngineDaemon_CP_1640_elements(22) & ReceiveEngineDaemon_CP_1640_elements(30) & ReceiveEngineDaemon_CP_1640_elements(45);
      gj_ReceiveEngineDaemon_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1640_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1052_update_start_
      -- CP-element group 44: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1052_Update/$entry
      -- CP-element group 44: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1052_Update/ccr
      -- 
    ccr_1864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(44), ack => call_stmt_1052_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1640_elements(46);
      gj_ReceiveEngineDaemon_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1640_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: marked-successors 
    -- CP-element group 45: 	40 
    -- CP-element group 45: 	43 
    -- CP-element group 45: 	20 
    -- CP-element group 45: 	28 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1052_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1052_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1052_Sample/cra
      -- 
    cra_1860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1052_call_ack_0, ack => ReceiveEngineDaemon_CP_1640_elements(45)); -- 
    -- CP-element group 46:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	11 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: 	16 
    -- CP-element group 46: 	15 
    -- CP-element group 46:  members (4) 
      -- CP-element group 46: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/$exit
      -- CP-element group 46: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1052_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1052_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/call_stmt_1052_Update/cca
      -- 
    cca_1865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1052_call_ack_1, ack => ReceiveEngineDaemon_CP_1640_elements(46)); -- 
    -- CP-element group 47:  transition  output  delay-element  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	14 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	10 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/condition_evaluated
      -- CP-element group 47: 	 branch_block_stmt_968/do_while_stmt_979/do_while_stmt_979_loop_body/loop_body_delay_to_condition_start
      -- 
    condition_evaluated_1752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(47), ack => do_while_stmt_979_branch_req_0); -- 
    -- Element group ReceiveEngineDaemon_CP_1640_elements(47) is a control-delay.
    cp_element_47_delay: control_delay_element  generic map(name => " 47_delay", delay_value => 1)  port map(req => ReceiveEngineDaemon_CP_1640_elements(14), ack => ReceiveEngineDaemon_CP_1640_elements(47), clk => clk, reset =>reset);
    -- CP-element group 48:  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	10 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_968/do_while_stmt_979/loop_exit/$exit
      -- CP-element group 48: 	 branch_block_stmt_968/do_while_stmt_979/loop_exit/ack
      -- 
    ack_1870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_979_branch_ack_0, ack => ReceiveEngineDaemon_CP_1640_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	10 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_968/do_while_stmt_979/loop_taken/$exit
      -- CP-element group 49: 	 branch_block_stmt_968/do_while_stmt_979/loop_taken/ack
      -- 
    ack_1874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_979_branch_ack_1, ack => ReceiveEngineDaemon_CP_1640_elements(49)); -- 
    -- CP-element group 50:  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	8 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	4 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_968/do_while_stmt_979/$exit
      -- 
    ReceiveEngineDaemon_CP_1640_elements(50) <= ReceiveEngineDaemon_CP_1640_elements(8);
    -- CP-element group 51:  merge  branch  transition  place  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	4 
    -- CP-element group 51: 	5 
    -- CP-element group 51: 	2 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	6 
    -- CP-element group 51: 	5 
    -- CP-element group 51:  members (49) 
      -- CP-element group 51: 	 branch_block_stmt_968/merge_stmt_970__exit__
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971__entry__
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_dead_link/$entry
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/$entry
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/$exit
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/$entry
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/$exit
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/$entry
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/$exit
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/BITSEL_u32_u1_974_inputs/$entry
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/BITSEL_u32_u1_974_inputs/$exit
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/BITSEL_u32_u1_974_inputs/RPIPE_CONTROL_REGISTER_972/$entry
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/BITSEL_u32_u1_974_inputs/RPIPE_CONTROL_REGISTER_972/$exit
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/BITSEL_u32_u1_974_inputs/RPIPE_CONTROL_REGISTER_972/Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/BITSEL_u32_u1_974_inputs/RPIPE_CONTROL_REGISTER_972/Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/BITSEL_u32_u1_974_inputs/RPIPE_CONTROL_REGISTER_972/Sample/req
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/BITSEL_u32_u1_974_inputs/RPIPE_CONTROL_REGISTER_972/Sample/ack
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/BITSEL_u32_u1_974_inputs/RPIPE_CONTROL_REGISTER_972/Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/BITSEL_u32_u1_974_inputs/RPIPE_CONTROL_REGISTER_972/Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/BITSEL_u32_u1_974_inputs/RPIPE_CONTROL_REGISTER_972/Update/req
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/BITSEL_u32_u1_974_inputs/RPIPE_CONTROL_REGISTER_972/Update/ack
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/SplitProtocol/$entry
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/SplitProtocol/$exit
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/SplitProtocol/Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/SplitProtocol/Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/SplitProtocol/Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/SplitProtocol/Sample/ra
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/SplitProtocol/Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/SplitProtocol/Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/SplitProtocol/Update/cr
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/BITSEL_u32_u1_974/SplitProtocol/Update/ca
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/SplitProtocol/$entry
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/SplitProtocol/$exit
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/SplitProtocol/Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/SplitProtocol/Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/SplitProtocol/Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/SplitProtocol/Sample/ra
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/SplitProtocol/Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/SplitProtocol/Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/SplitProtocol/Update/cr
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/NOT_u1_u1_975/SplitProtocol/Update/ca
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_eval_test/branch_req
      -- CP-element group 51: 	 branch_block_stmt_968/NOT_u1_u1_975_place
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_if_link/$entry
      -- CP-element group 51: 	 branch_block_stmt_968/if_stmt_971_else_link/$entry
      -- CP-element group 51: 	 branch_block_stmt_968/merge_stmt_970_PhiReqMerge
      -- CP-element group 51: 	 branch_block_stmt_968/merge_stmt_970_PhiAck/$entry
      -- CP-element group 51: 	 branch_block_stmt_968/merge_stmt_970_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_968/merge_stmt_970_PhiAck/dummy
      -- 
    branch_req_1727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1640_elements(51), ack => if_stmt_971_branch_req_0); -- 
    ReceiveEngineDaemon_CP_1640_elements(51) <= OrReduce(ReceiveEngineDaemon_CP_1640_elements(4) & ReceiveEngineDaemon_CP_1640_elements(5) & ReceiveEngineDaemon_CP_1640_elements(2));
    ReceiveEngineDaemon_do_while_stmt_979_terminator_1875: loop_terminator -- 
      generic map (name => " ReceiveEngineDaemon_do_while_stmt_979_terminator_1875", max_iterations_in_flight =>31) 
      port map(loop_body_exit => ReceiveEngineDaemon_CP_1640_elements(11),loop_continue => ReceiveEngineDaemon_CP_1640_elements(49),loop_terminate => ReceiveEngineDaemon_CP_1640_elements(48),loop_back => ReceiveEngineDaemon_CP_1640_elements(9),loop_exit => ReceiveEngineDaemon_CP_1640_elements(8),clk => clk, reset => reset); -- 
    entry_tmerge_1753_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= ReceiveEngineDaemon_CP_1640_elements(12);
        preds(1)  <= ReceiveEngineDaemon_CP_1640_elements(13);
        entry_tmerge_1753 : transition_merge -- 
          generic map(name => " entry_tmerge_1753")
          port map (preds => preds, symbol_out => ReceiveEngineDaemon_CP_1640_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_1057_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_974_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1002_1002_delayed_10_0_1019 : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1013_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_975_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_995_995_delayed_10_0_1009 : std_logic_vector(0 downto 0);
    signal RPIPE_CONTROL_REGISTER_1055_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CONTROL_REGISTER_972_wire : std_logic_vector(31 downto 0);
    signal RPIPE_FREE_Q_1048_wire : std_logic_vector(35 downto 0);
    signal RPIPE_FREE_Q_984_wire : std_logic_vector(35 downto 0);
    signal bad_packet_identifier_1005 : std_logic_vector(0 downto 0);
    signal cond_1029 : std_logic_vector(0 downto 0);
    signal free_flag_1024 : std_logic_vector(0 downto 0);
    signal konst_1027_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1056_wire_constant : std_logic_vector(31 downto 0);
    signal konst_966_wire_constant : std_logic_vector(5 downto 0);
    signal konst_973_wire_constant : std_logic_vector(31 downto 0);
    signal ok_flag_1015 : std_logic_vector(0 downto 0);
    signal push_status_1052 : std_logic_vector(0 downto 0);
    signal rx_buffer_pointer_32_987 : std_logic_vector(31 downto 0);
    signal rx_buffer_pointer_36_1016_delayed_10_0_1036 : std_logic_vector(35 downto 0);
    signal rx_buffer_pointer_36_1024_delayed_10_0_1044 : std_logic_vector(35 downto 0);
    signal rx_buffer_pointer_36_995 : std_logic_vector(35 downto 0);
    signal slice_1050_wire : std_logic_vector(31 downto 0);
    signal status_987 : std_logic_vector(0 downto 0);
    signal type_cast_1047_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_983_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_993_wire_constant : std_logic_vector(3 downto 0);
    -- 
  begin -- 
    konst_1027_wire_constant <= "1";
    konst_1056_wire_constant <= "00000000000000000000000000000000";
    konst_966_wire_constant <= "000000";
    konst_973_wire_constant <= "00000000000000000000000000000000";
    type_cast_1047_wire_constant <= "1";
    type_cast_983_wire_constant <= "1";
    type_cast_993_wire_constant <= "0000";
    -- flow-through slice operator slice_1050_inst
    slice_1050_wire <= rx_buffer_pointer_36_1024_delayed_10_0_1044(35 downto 4);
    W_rx_buffer_pointer_36_1016_delayed_10_0_1034_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_36_1016_delayed_10_0_1034_inst_req_0;
      W_rx_buffer_pointer_36_1016_delayed_10_0_1034_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_36_1016_delayed_10_0_1034_inst_req_1;
      W_rx_buffer_pointer_36_1016_delayed_10_0_1034_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_36_1016_delayed_10_0_1034_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_36_1016_delayed_10_0_1034_inst",
        buffer_size => 10,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_36_995,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_36_1016_delayed_10_0_1036,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_36_1024_delayed_10_0_1042_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_36_1024_delayed_10_0_1042_inst_req_0;
      W_rx_buffer_pointer_36_1024_delayed_10_0_1042_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_36_1024_delayed_10_0_1042_inst_req_1;
      W_rx_buffer_pointer_36_1024_delayed_10_0_1042_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_36_1024_delayed_10_0_1042_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_36_1024_delayed_10_0_1042_inst",
        buffer_size => 10,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_36_995,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_36_1024_delayed_10_0_1044,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_979_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_1057_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_979_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_979_branch_req_0,
          ack0 => do_while_stmt_979_branch_ack_0,
          ack1 => do_while_stmt_979_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_971_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_975_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_971_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_971_branch_req_0,
          ack0 => if_stmt_971_branch_ack_0,
          ack1 => if_stmt_971_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_1014_inst
    process(NOT_u1_u1_995_995_delayed_10_0_1009, NOT_u1_u1_1013_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_995_995_delayed_10_0_1009, NOT_u1_u1_1013_wire, tmp_var);
      ok_flag_1015 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1023_inst
    process(NOT_u1_u1_1002_1002_delayed_10_0_1019, bad_packet_identifier_1005) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_1002_1002_delayed_10_0_1019, bad_packet_identifier_1005, tmp_var);
      free_flag_1024 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1057_inst
    process(RPIPE_CONTROL_REGISTER_1055_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1055_wire, konst_1056_wire_constant, tmp_var);
      BITSEL_u32_u1_1057_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_974_inst
    process(RPIPE_CONTROL_REGISTER_972_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_972_wire, konst_973_wire_constant, tmp_var);
      BITSEL_u32_u1_974_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u36_994_inst
    process(rx_buffer_pointer_32_987) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(rx_buffer_pointer_32_987, type_cast_993_wire_constant, tmp_var);
      rx_buffer_pointer_36_995 <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1028_inst
    process(ok_flag_1015) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ok_flag_1015, konst_1027_wire_constant, tmp_var);
      cond_1029 <= tmp_var; --
    end process;
    -- shared split operator group (6) : NOT_u1_u1_1008_inst 
    ApIntNot_group_6: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 10);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= status_987;
      NOT_u1_u1_995_995_delayed_10_0_1009 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1008_inst_req_0;
      NOT_u1_u1_1008_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1008_inst_req_1;
      NOT_u1_u1_1008_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_6_gI: SplitGuardInterface generic map(name => "ApIntNot_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 10,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- unary operator NOT_u1_u1_1013_inst
    process(bad_packet_identifier_1005) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", bad_packet_identifier_1005, tmp_var);
      NOT_u1_u1_1013_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (8) : NOT_u1_u1_1018_inst 
    ApIntNot_group_8: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 10);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= status_987;
      NOT_u1_u1_1002_1002_delayed_10_0_1019 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1018_inst_req_0;
      NOT_u1_u1_1018_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1018_inst_req_1;
      NOT_u1_u1_1018_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_8_gI: SplitGuardInterface generic map(name => "ApIntNot_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 10,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- unary operator NOT_u1_u1_975_inst
    process(BITSEL_u32_u1_974_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_974_wire, tmp_var);
      NOT_u1_u1_975_wire <= tmp_var; -- 
    end process;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1055_wire <= CONTROL_REGISTER;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_972_wire <= CONTROL_REGISTER;
    -- read from input-signal FREE_Q
    RPIPE_FREE_Q_1048_wire <= FREE_Q;
    RPIPE_FREE_Q_984_wire <= FREE_Q;
    -- shared outport operator group (0) : WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_inst_req_0;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_inst_req_1;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_965_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_966_wire_constant;
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_WRITTEN_RX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(5 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1005_call 
    loadBuffer_call_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 10);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1005_call_req_0;
      call_stmt_1005_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1005_call_req_1;
      call_stmt_1005_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not status_987(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadBuffer_call_group_0_gI: SplitGuardInterface generic map(name => "loadBuffer_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_36_995;
      bad_packet_identifier_1005 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadBuffer_call_reqs(0),
          ackR => loadBuffer_call_acks(0),
          dataR => loadBuffer_call_data(35 downto 0),
          tagR => loadBuffer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => loadBuffer_return_acks(0), -- cross-over
          ackL => loadBuffer_return_reqs(0), -- cross-over
          dataL => loadBuffer_return_data(0 downto 0),
          tagL => loadBuffer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1039_call 
    populateRxQueue_call_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1039_call_req_0;
      call_stmt_1039_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1039_call_req_1;
      call_stmt_1039_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ok_flag_1015(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      populateRxQueue_call_group_1_gI: SplitGuardInterface generic map(name => "populateRxQueue_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_36_1016_delayed_10_0_1036;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => populateRxQueue_call_reqs(0),
          ackR => populateRxQueue_call_acks(0),
          dataR => populateRxQueue_call_data(35 downto 0),
          tagR => populateRxQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => populateRxQueue_return_acks(0), -- cross-over
          ackL => populateRxQueue_return_reqs(0), -- cross-over
          tagL => populateRxQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1052_call 
    pushIntoQueue_call_group_2: Block -- 
      signal data_in: std_logic_vector(68 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1052_call_req_0;
      call_stmt_1052_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1052_call_req_1;
      call_stmt_1052_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= free_flag_1024(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_2_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1047_wire_constant & RPIPE_FREE_Q_1048_wire & slice_1050_wire;
      push_status_1052 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 69,
        owidth => 69,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(68 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_987_call 
    popFromQueue_call_group_3: Block -- 
      signal data_in: std_logic_vector(36 downto 0);
      signal data_out: std_logic_vector(32 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_987_call_req_0;
      call_stmt_987_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_987_call_req_1;
      call_stmt_987_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      popFromQueue_call_group_3_gI: SplitGuardInterface generic map(name => "popFromQueue_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_983_wire_constant & RPIPE_FREE_Q_984_wire;
      rx_buffer_pointer_32_987 <= data_out(32 downto 1);
      status_987 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 37,
        owidth => 37,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => popFromQueue_call_reqs(0),
          ackR => popFromQueue_call_acks(0),
          dataR => popFromQueue_call_data(36 downto 0),
          tagR => popFromQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 33,
          owidth => 33,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => popFromQueue_return_acks(0), -- cross-over
          ackL => popFromQueue_return_reqs(0), -- cross-over
          dataL => popFromQueue_return_data(32 downto 0),
          tagL => popFromQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end ReceiveEngineDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity SoftwareRegisterAccessDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    AFB_NIC_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_read_data : in   std_logic_vector(73 downto 0);
    FREE_Q_pipe_write_req : out  std_logic_vector(0 downto 0);
    FREE_Q_pipe_write_ack : in   std_logic_vector(0 downto 0);
    FREE_Q_pipe_write_data : out  std_logic_vector(35 downto 0);
    AFB_NIC_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_write_data : out  std_logic_vector(32 downto 0);
    CONTROL_REGISTER_pipe_write_req : out  std_logic_vector(0 downto 0);
    CONTROL_REGISTER_pipe_write_ack : in   std_logic_vector(0 downto 0);
    CONTROL_REGISTER_pipe_write_data : out  std_logic_vector(31 downto 0);
    NUMBER_OF_SERVERS_pipe_write_req : out  std_logic_vector(0 downto 0);
    NUMBER_OF_SERVERS_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NUMBER_OF_SERVERS_pipe_write_data : out  std_logic_vector(31 downto 0);
    UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
    UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
    UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
    UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity SoftwareRegisterAccessDaemon;
architecture SoftwareRegisterAccessDaemon_arch of SoftwareRegisterAccessDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal SoftwareRegisterAccessDaemon_CP_1894_start: Boolean;
  signal SoftwareRegisterAccessDaemon_CP_1894_symbol: Boolean;
  -- volatile/operator module components. 
  component UpdateRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      bmask : in  std_logic_vector(3 downto 0);
      rval : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      index : in  std_logic_vector(5 downto 0);
      wval : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal phi_stmt_1082_ack_0 : boolean;
  signal phi_stmt_1072_req_1 : boolean;
  signal check_num_server_1196_1086_buf_ack_0 : boolean;
  signal check_num_server_1196_1086_buf_ack_1 : boolean;
  signal phi_stmt_1066_req_0 : boolean;
  signal phi_stmt_1066_req_1 : boolean;
  signal do_while_stmt_1064_branch_req_0 : boolean;
  signal phi_stmt_1066_ack_0 : boolean;
  signal array_obj_ref_1122_load_0_req_1 : boolean;
  signal array_obj_ref_1091_load_0_req_0 : boolean;
  signal check_num_server_1196_1086_buf_req_1 : boolean;
  signal array_obj_ref_1122_load_0_ack_1 : boolean;
  signal array_obj_ref_1122_load_0_req_0 : boolean;
  signal array_obj_ref_1122_load_0_ack_0 : boolean;
  signal check_control_regsiter_1178_1076_buf_ack_0 : boolean;
  signal check_control_regsiter_1178_1076_buf_req_0 : boolean;
  signal check_num_server_1196_1086_buf_req_0 : boolean;
  signal phi_stmt_1082_req_1 : boolean;
  signal phi_stmt_1077_ack_0 : boolean;
  signal check_free_q_1187_1081_buf_ack_1 : boolean;
  signal phi_stmt_1077_req_1 : boolean;
  signal check_free_q_1187_1081_buf_req_1 : boolean;
  signal phi_stmt_1082_req_0 : boolean;
  signal phi_stmt_1077_req_0 : boolean;
  signal array_obj_ref_1091_load_0_ack_1 : boolean;
  signal phi_stmt_1072_ack_0 : boolean;
  signal check_free_q_1187_1081_buf_ack_0 : boolean;
  signal array_obj_ref_1091_load_0_req_1 : boolean;
  signal check_control_regsiter_1178_1076_buf_ack_1 : boolean;
  signal check_control_regsiter_1178_1076_buf_req_1 : boolean;
  signal phi_stmt_1072_req_0 : boolean;
  signal check_free_q_1187_1081_buf_req_0 : boolean;
  signal array_obj_ref_1091_load_0_ack_0 : boolean;
  signal WPIPE_CONTROL_REGISTER_1120_inst_req_0 : boolean;
  signal WPIPE_CONTROL_REGISTER_1120_inst_ack_0 : boolean;
  signal WPIPE_CONTROL_REGISTER_1120_inst_req_1 : boolean;
  signal WPIPE_CONTROL_REGISTER_1120_inst_ack_1 : boolean;
  signal array_obj_ref_1127_load_0_req_0 : boolean;
  signal array_obj_ref_1127_load_0_ack_0 : boolean;
  signal array_obj_ref_1127_load_0_req_1 : boolean;
  signal array_obj_ref_1127_load_0_ack_1 : boolean;
  signal W_update_free_q_pipe_1104_delayed_5_0_1129_inst_req_0 : boolean;
  signal W_update_free_q_pipe_1104_delayed_5_0_1129_inst_ack_0 : boolean;
  signal W_update_free_q_pipe_1104_delayed_5_0_1129_inst_req_1 : boolean;
  signal W_update_free_q_pipe_1104_delayed_5_0_1129_inst_ack_1 : boolean;
  signal type_cast_1138_inst_req_0 : boolean;
  signal type_cast_1138_inst_ack_0 : boolean;
  signal type_cast_1138_inst_req_1 : boolean;
  signal type_cast_1138_inst_ack_1 : boolean;
  signal WPIPE_FREE_Q_1133_inst_req_0 : boolean;
  signal WPIPE_FREE_Q_1133_inst_ack_0 : boolean;
  signal WPIPE_FREE_Q_1133_inst_req_1 : boolean;
  signal WPIPE_FREE_Q_1133_inst_ack_1 : boolean;
  signal array_obj_ref_1143_load_0_req_0 : boolean;
  signal array_obj_ref_1143_load_0_ack_0 : boolean;
  signal array_obj_ref_1143_load_0_req_1 : boolean;
  signal array_obj_ref_1143_load_0_ack_1 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1141_inst_req_0 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1141_inst_ack_0 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1141_inst_req_1 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1141_inst_ack_1 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1146_inst_req_0 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1146_inst_ack_0 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1146_inst_req_1 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1146_inst_ack_1 : boolean;
  signal array_obj_ref_1199_load_0_req_0 : boolean;
  signal array_obj_ref_1199_load_0_ack_0 : boolean;
  signal array_obj_ref_1199_load_0_req_1 : boolean;
  signal array_obj_ref_1199_load_0_ack_1 : boolean;
  signal W_rwbar_1177_delayed_5_0_1201_inst_req_0 : boolean;
  signal W_rwbar_1177_delayed_5_0_1201_inst_ack_0 : boolean;
  signal W_rwbar_1177_delayed_5_0_1201_inst_req_1 : boolean;
  signal W_rwbar_1177_delayed_5_0_1201_inst_ack_1 : boolean;
  signal W_bmask_1178_delayed_5_0_1204_inst_req_0 : boolean;
  signal W_bmask_1178_delayed_5_0_1204_inst_ack_0 : boolean;
  signal W_bmask_1178_delayed_5_0_1204_inst_req_1 : boolean;
  signal W_bmask_1178_delayed_5_0_1204_inst_ack_1 : boolean;
  signal W_wdata_1180_delayed_5_0_1207_inst_req_0 : boolean;
  signal W_wdata_1180_delayed_5_0_1207_inst_ack_0 : boolean;
  signal W_wdata_1180_delayed_5_0_1207_inst_req_1 : boolean;
  signal W_wdata_1180_delayed_5_0_1207_inst_ack_1 : boolean;
  signal W_index_1181_delayed_5_0_1210_inst_req_0 : boolean;
  signal W_index_1181_delayed_5_0_1210_inst_ack_0 : boolean;
  signal W_index_1181_delayed_5_0_1210_inst_req_1 : boolean;
  signal W_index_1181_delayed_5_0_1210_inst_ack_1 : boolean;
  signal call_stmt_1219_call_req_0 : boolean;
  signal call_stmt_1219_call_ack_0 : boolean;
  signal call_stmt_1219_call_req_1 : boolean;
  signal call_stmt_1219_call_ack_1 : boolean;
  signal W_rwbar_1185_delayed_5_0_1220_inst_req_0 : boolean;
  signal W_rwbar_1185_delayed_5_0_1220_inst_ack_0 : boolean;
  signal W_rwbar_1185_delayed_5_0_1220_inst_req_1 : boolean;
  signal W_rwbar_1185_delayed_5_0_1220_inst_ack_1 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1236_inst_req_0 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1236_inst_ack_0 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1236_inst_req_1 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1236_inst_ack_1 : boolean;
  signal do_while_stmt_1064_branch_ack_0 : boolean;
  signal do_while_stmt_1064_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "SoftwareRegisterAccessDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  SoftwareRegisterAccessDaemon_CP_1894_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "SoftwareRegisterAccessDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= SoftwareRegisterAccessDaemon_CP_1894_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= SoftwareRegisterAccessDaemon_CP_1894_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= SoftwareRegisterAccessDaemon_CP_1894_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  SoftwareRegisterAccessDaemon_CP_1894: Block -- control-path 
    signal SoftwareRegisterAccessDaemon_CP_1894_elements: BooleanArray(166 downto 0);
    -- 
  begin -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(0) <= SoftwareRegisterAccessDaemon_CP_1894_start;
    SoftwareRegisterAccessDaemon_CP_1894_symbol <= SoftwareRegisterAccessDaemon_CP_1894_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1063/do_while_stmt_1064__entry__
      -- CP-element group 0: 	 branch_block_stmt_1063/$entry
      -- CP-element group 0: 	 branch_block_stmt_1063/branch_block_stmt_1063__entry__
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	166 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1063/do_while_stmt_1064__exit__
      -- CP-element group 1: 	 branch_block_stmt_1063/$exit
      -- CP-element group 1: 	 branch_block_stmt_1063/branch_block_stmt_1063__exit__
      -- CP-element group 1: 	 $exit
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(1) <= SoftwareRegisterAccessDaemon_CP_1894_elements(166);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064__entry__
      -- CP-element group 2: 	 branch_block_stmt_1063/do_while_stmt_1064/$entry
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(2) <= SoftwareRegisterAccessDaemon_CP_1894_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	166 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064__exit__
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1063/do_while_stmt_1064/loop_back
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	164 
    -- CP-element group 5: 	165 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1063/do_while_stmt_1064/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1063/do_while_stmt_1064/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1063/do_while_stmt_1064/loop_taken/$entry
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(5) <= SoftwareRegisterAccessDaemon_CP_1894_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	163 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1063/do_while_stmt_1064/loop_body_done
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(6) <= SoftwareRegisterAccessDaemon_CP_1894_elements(163);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	38 
    -- CP-element group 7: 	57 
    -- CP-element group 7: 	76 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/back_edge_to_loop_body
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(7) <= SoftwareRegisterAccessDaemon_CP_1894_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	40 
    -- CP-element group 8: 	59 
    -- CP-element group 8: 	78 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/first_time_through_loop_body
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(8) <= SoftwareRegisterAccessDaemon_CP_1894_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	33 
    -- CP-element group 9: 	122 
    -- CP-element group 9: 	157 
    -- CP-element group 9: 	115 
    -- CP-element group 9: 	93 
    -- CP-element group 9: 	100 
    -- CP-element group 9: 	51 
    -- CP-element group 9: 	52 
    -- CP-element group 9: 	70 
    -- CP-element group 9: 	71 
    -- CP-element group 9: 	89 
    -- CP-element group 9:  members (10) 
      -- CP-element group 9: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_root_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_root_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_root_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_root_address_calculated
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	157 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/condition_evaluated
      -- 
    condition_evaluated_1918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(10), ack => do_while_stmt_1064_branch_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(14) & SoftwareRegisterAccessDaemon_CP_1894_elements(157);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	32 
    -- CP-element group 11: 	51 
    -- CP-element group 11: 	70 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	72 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1066_sample_start__ps
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 31,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(15) & SoftwareRegisterAccessDaemon_CP_1894_elements(32) & SoftwareRegisterAccessDaemon_CP_1894_elements(51) & SoftwareRegisterAccessDaemon_CP_1894_elements(70) & SoftwareRegisterAccessDaemon_CP_1894_elements(14);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	54 
    -- CP-element group 12: 	73 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	123 
    -- CP-element group 12: 	163 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	32 
    -- CP-element group 12: 	51 
    -- CP-element group 12: 	70 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1077_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1066_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1072_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1082_sample_completed_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(17) & SoftwareRegisterAccessDaemon_CP_1894_elements(35) & SoftwareRegisterAccessDaemon_CP_1894_elements(54) & SoftwareRegisterAccessDaemon_CP_1894_elements(73);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	33 
    -- CP-element group 13: 	52 
    -- CP-element group 13: 	71 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	36 
    -- CP-element group 13: 	55 
    -- CP-element group 13: 	74 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1066_update_start__ps
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(16) & SoftwareRegisterAccessDaemon_CP_1894_elements(33) & SoftwareRegisterAccessDaemon_CP_1894_elements(52) & SoftwareRegisterAccessDaemon_CP_1894_elements(71);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	56 
    -- CP-element group 14: 	75 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/aggregated_phi_update_ack
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(18) & SoftwareRegisterAccessDaemon_CP_1894_elements(37) & SoftwareRegisterAccessDaemon_CP_1894_elements(56) & SoftwareRegisterAccessDaemon_CP_1894_elements(75);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1066_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(9) & SoftwareRegisterAccessDaemon_CP_1894_elements(12);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	120 
    -- CP-element group 16: 	117 
    -- CP-element group 16: 	102 
    -- CP-element group 16: 	106 
    -- CP-element group 16: 	98 
    -- CP-element group 16: 	95 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1066_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(9) & SoftwareRegisterAccessDaemon_CP_1894_elements(120) & SoftwareRegisterAccessDaemon_CP_1894_elements(117) & SoftwareRegisterAccessDaemon_CP_1894_elements(102) & SoftwareRegisterAccessDaemon_CP_1894_elements(106) & SoftwareRegisterAccessDaemon_CP_1894_elements(98) & SoftwareRegisterAccessDaemon_CP_1894_elements(95);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1066_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	119 
    -- CP-element group 18: 	115 
    -- CP-element group 18: 	93 
    -- CP-element group 18: 	104 
    -- CP-element group 18: 	97 
    -- CP-element group 18: 	100 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1066_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1066_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1066_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(19) <= SoftwareRegisterAccessDaemon_CP_1894_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1066_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1066_loopback_sample_req_ps
      -- 
    phi_stmt_1066_loopback_sample_req_1933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1066_loopback_sample_req_1933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(20), ack => phi_stmt_1066_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1066_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(21) <= SoftwareRegisterAccessDaemon_CP_1894_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1066_entry_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1066_entry_sample_req
      -- 
    phi_stmt_1066_entry_sample_req_1936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1066_entry_sample_req_1936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(22), ack => phi_stmt_1066_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1066_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1066_phi_mux_ack_ps
      -- 
    phi_stmt_1066_phi_mux_ack_1939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1066_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1069_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1069_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1069_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1069_sample_start_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1069_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1069_update_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1069_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(26) <= SoftwareRegisterAccessDaemon_CP_1894_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1069_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1894_elements(25), ack => SoftwareRegisterAccessDaemon_CP_1894_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1071_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1071_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1071_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1071_sample_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1071_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1071_update_start_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1071_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(30) <= SoftwareRegisterAccessDaemon_CP_1894_elements(31);
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	30 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1071_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1894_elements(29), ack => SoftwareRegisterAccessDaemon_CP_1894_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	12 
    -- CP-element group 32: 	125 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	11 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1072_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(9) & SoftwareRegisterAccessDaemon_CP_1894_elements(12) & SoftwareRegisterAccessDaemon_CP_1894_elements(125);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	9 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	98 
    -- CP-element group 33: 	95 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1072_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(9) & SoftwareRegisterAccessDaemon_CP_1894_elements(98) & SoftwareRegisterAccessDaemon_CP_1894_elements(95);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1072_sample_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(34) <= SoftwareRegisterAccessDaemon_CP_1894_elements(11);
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1072_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(35) is bound as output of CP function.
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	13 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1072_update_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(36) <= SoftwareRegisterAccessDaemon_CP_1894_elements(13);
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: 	93 
    -- CP-element group 37: 	97 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1072_update_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1072_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	7 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1072_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(38) <= SoftwareRegisterAccessDaemon_CP_1894_elements(7);
    -- CP-element group 39:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1072_loopback_sample_req
      -- CP-element group 39: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1072_loopback_sample_req_ps
      -- 
    phi_stmt_1072_loopback_sample_req_1967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1072_loopback_sample_req_1967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(39), ack => phi_stmt_1072_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	8 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1072_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(40) <= SoftwareRegisterAccessDaemon_CP_1894_elements(8);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1072_entry_sample_req_ps
      -- CP-element group 41: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1072_entry_sample_req
      -- 
    phi_stmt_1072_entry_sample_req_1970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1072_entry_sample_req_1970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(41), ack => phi_stmt_1072_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1072_phi_mux_ack_ps
      -- CP-element group 42: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1072_phi_mux_ack
      -- 
    phi_stmt_1072_phi_mux_ack_1973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1072_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1075_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1075_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1075_sample_completed__ps
      -- CP-element group 43: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1075_sample_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1075_update_start_
      -- CP-element group 44: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1075_update_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1075_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(45) <= SoftwareRegisterAccessDaemon_CP_1894_elements(46);
    -- CP-element group 46:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	45 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1075_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(46) is a control-delay.
    cp_element_46_delay: control_delay_element  generic map(name => " 46_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1894_elements(44), ack => SoftwareRegisterAccessDaemon_CP_1894_elements(46), clk => clk, reset =>reset);
    -- CP-element group 47:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_control_regsiter_1076_Sample/req
      -- CP-element group 47: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_control_regsiter_1076_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_control_regsiter_1076_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_control_regsiter_1076_sample_start__ps
      -- 
    req_1994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(47), ack => check_control_regsiter_1178_1076_buf_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_control_regsiter_1076_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_control_regsiter_1076_update_start_
      -- CP-element group 48: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_control_regsiter_1076_update_start__ps
      -- CP-element group 48: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_control_regsiter_1076_Update/req
      -- 
    req_1999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(48), ack => check_control_regsiter_1178_1076_buf_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_control_regsiter_1076_Sample/ack
      -- CP-element group 49: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_control_regsiter_1076_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_control_regsiter_1076_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_control_regsiter_1076_sample_completed__ps
      -- 
    ack_1995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_control_regsiter_1178_1076_buf_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(49)); -- 
    -- CP-element group 50:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_control_regsiter_1076_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_control_regsiter_1076_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_control_regsiter_1076_update_completed__ps
      -- CP-element group 50: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_control_regsiter_1076_Update/ack
      -- 
    ack_2000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_control_regsiter_1178_1076_buf_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(50)); -- 
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	9 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	12 
    -- CP-element group 51: 	125 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	11 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1077_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(9) & SoftwareRegisterAccessDaemon_CP_1894_elements(12) & SoftwareRegisterAccessDaemon_CP_1894_elements(125);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	9 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	102 
    -- CP-element group 52: 	106 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	13 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1077_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(9) & SoftwareRegisterAccessDaemon_CP_1894_elements(102) & SoftwareRegisterAccessDaemon_CP_1894_elements(106);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	11 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1077_sample_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(53) <= SoftwareRegisterAccessDaemon_CP_1894_elements(11);
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	12 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1077_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(54) is bound as output of CP function.
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	13 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1077_update_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(55) <= SoftwareRegisterAccessDaemon_CP_1894_elements(13);
    -- CP-element group 56:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	14 
    -- CP-element group 56: 	104 
    -- CP-element group 56: 	100 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1077_update_completed__ps
      -- CP-element group 56: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1077_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	7 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1077_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(57) <= SoftwareRegisterAccessDaemon_CP_1894_elements(7);
    -- CP-element group 58:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1077_loopback_sample_req_ps
      -- CP-element group 58: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1077_loopback_sample_req
      -- 
    phi_stmt_1077_loopback_sample_req_2011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1077_loopback_sample_req_2011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(58), ack => phi_stmt_1077_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	8 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1077_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(59) <= SoftwareRegisterAccessDaemon_CP_1894_elements(8);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1077_entry_sample_req_ps
      -- CP-element group 60: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1077_entry_sample_req
      -- 
    phi_stmt_1077_entry_sample_req_2014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1077_entry_sample_req_2014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(60), ack => phi_stmt_1077_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1077_phi_mux_ack_ps
      -- CP-element group 61: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1077_phi_mux_ack
      -- 
    phi_stmt_1077_phi_mux_ack_2017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1077_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1080_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1080_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1080_sample_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1080_sample_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1080_update_start__ps
      -- CP-element group 63: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1080_update_start_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1080_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(64) <= SoftwareRegisterAccessDaemon_CP_1894_elements(65);
    -- CP-element group 65:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	64 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1080_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(65) is a control-delay.
    cp_element_65_delay: control_delay_element  generic map(name => " 65_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1894_elements(63), ack => SoftwareRegisterAccessDaemon_CP_1894_elements(65), clk => clk, reset =>reset);
    -- CP-element group 66:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_free_q_1081_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_free_q_1081_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_free_q_1081_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_free_q_1081_Sample/req
      -- 
    req_2038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(66), ack => check_free_q_1187_1081_buf_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_free_q_1081_update_start_
      -- CP-element group 67: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_free_q_1081_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_free_q_1081_Update/req
      -- CP-element group 67: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_free_q_1081_Update/$entry
      -- 
    req_2043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(67), ack => check_free_q_1187_1081_buf_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_free_q_1081_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_free_q_1081_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_free_q_1081_Sample/ack
      -- CP-element group 68: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_free_q_1081_Sample/$exit
      -- 
    ack_2039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_free_q_1187_1081_buf_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(68)); -- 
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_free_q_1081_update_completed__ps
      -- CP-element group 69: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_free_q_1081_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_free_q_1081_Update/ack
      -- CP-element group 69: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_free_q_1081_Update/$exit
      -- 
    ack_2044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_free_q_1187_1081_buf_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(69)); -- 
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	9 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	12 
    -- CP-element group 70: 	125 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	11 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1082_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(9) & SoftwareRegisterAccessDaemon_CP_1894_elements(12) & SoftwareRegisterAccessDaemon_CP_1894_elements(125);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	9 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	120 
    -- CP-element group 71: 	117 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	13 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1082_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(9) & SoftwareRegisterAccessDaemon_CP_1894_elements(120) & SoftwareRegisterAccessDaemon_CP_1894_elements(117);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	11 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1082_sample_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(72) <= SoftwareRegisterAccessDaemon_CP_1894_elements(11);
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	12 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1082_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(73) is bound as output of CP function.
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	13 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1082_update_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(74) <= SoftwareRegisterAccessDaemon_CP_1894_elements(13);
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	14 
    -- CP-element group 75: 	119 
    -- CP-element group 75: 	115 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1082_update_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1082_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	7 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1082_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(76) <= SoftwareRegisterAccessDaemon_CP_1894_elements(7);
    -- CP-element group 77:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1082_loopback_sample_req_ps
      -- CP-element group 77: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1082_loopback_sample_req
      -- 
    phi_stmt_1082_loopback_sample_req_2055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1082_loopback_sample_req_2055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(77), ack => phi_stmt_1082_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	8 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1082_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(78) <= SoftwareRegisterAccessDaemon_CP_1894_elements(8);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1082_entry_sample_req_ps
      -- CP-element group 79: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1082_entry_sample_req
      -- 
    phi_stmt_1082_entry_sample_req_2058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1082_entry_sample_req_2058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(79), ack => phi_stmt_1082_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(79) is bound as output of CP function.
    -- CP-element group 80:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1082_phi_mux_ack
      -- CP-element group 80: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/phi_stmt_1082_phi_mux_ack_ps
      -- 
    phi_stmt_1082_phi_mux_ack_2061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1082_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(80)); -- 
    -- CP-element group 81:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1085_sample_completed__ps
      -- CP-element group 81: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1085_sample_start__ps
      -- CP-element group 81: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1085_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1085_sample_start_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1085_update_start__ps
      -- CP-element group 82: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1085_update_start_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(82) is bound as output of CP function.
    -- CP-element group 83:  join  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1085_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(83) <= SoftwareRegisterAccessDaemon_CP_1894_elements(84);
    -- CP-element group 84:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	83 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1085_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1894_elements(82), ack => SoftwareRegisterAccessDaemon_CP_1894_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_num_server_1086_sample_start__ps
      -- CP-element group 85: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_num_server_1086_Sample/req
      -- CP-element group 85: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_num_server_1086_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_num_server_1086_sample_start_
      -- 
    req_2082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(85), ack => check_num_server_1196_1086_buf_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (4) 
      -- CP-element group 86: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_num_server_1086_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_num_server_1086_update_start__ps
      -- CP-element group 86: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_num_server_1086_Update/req
      -- CP-element group 86: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_num_server_1086_update_start_
      -- 
    req_2087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(86), ack => check_num_server_1196_1086_buf_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_num_server_1086_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_num_server_1086_sample_completed__ps
      -- CP-element group 87: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_num_server_1086_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_num_server_1086_sample_completed_
      -- 
    ack_2083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_num_server_1196_1086_buf_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(87)); -- 
    -- CP-element group 88:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_num_server_1086_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_num_server_1086_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_num_server_1086_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/R_check_num_server_1086_update_completed__ps
      -- 
    ack_2088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_num_server_1196_1086_buf_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	9 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: 	149 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Sample/word_access_start/word_0/rr
      -- CP-element group 89: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Sample/word_access_start/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Sample/word_access_start/$entry
      -- CP-element group 89: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Sample/$entry
      -- 
    rr_2106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(89), ack => array_obj_ref_1091_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(9) & SoftwareRegisterAccessDaemon_CP_1894_elements(91) & SoftwareRegisterAccessDaemon_CP_1894_elements(149);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_update_start_
      -- CP-element group 90: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Update/word_access_complete/word_0/$entry
      -- CP-element group 90: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Update/word_access_complete/$entry
      -- CP-element group 90: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Update/word_access_complete/word_0/cr
      -- 
    cr_2117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(90), ack => array_obj_ref_1091_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1894_elements(92);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	158 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Sample/word_access_start/word_0/$exit
      -- CP-element group 91: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Sample/word_access_start/$exit
      -- CP-element group 91: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Sample/word_access_start/word_0/ra
      -- 
    ra_2107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1091_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(91)); -- 
    -- CP-element group 92:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	163 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Update/array_obj_ref_1091_Merge/merge_req
      -- CP-element group 92: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Update/array_obj_ref_1091_Merge/$entry
      -- CP-element group 92: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Update/array_obj_ref_1091_Merge/merge_ack
      -- CP-element group 92: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Update/word_access_complete/$exit
      -- CP-element group 92: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Update/word_access_complete/word_0/$exit
      -- CP-element group 92: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Update/word_access_complete/word_0/ca
      -- CP-element group 92: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_Update/array_obj_ref_1091_Merge/$exit
      -- 
    ca_2118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1091_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	9 
    -- CP-element group 93: 	18 
    -- CP-element group 93: 	37 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	149 
    -- CP-element group 93: 	95 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Sample/word_access_start/word_0/rr
      -- CP-element group 93: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Sample/word_access_start/$entry
      -- CP-element group 93: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Sample/word_access_start/word_0/$entry
      -- 
    rr_2140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(93), ack => array_obj_ref_1122_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(9) & SoftwareRegisterAccessDaemon_CP_1894_elements(18) & SoftwareRegisterAccessDaemon_CP_1894_elements(37) & SoftwareRegisterAccessDaemon_CP_1894_elements(149) & SoftwareRegisterAccessDaemon_CP_1894_elements(95);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	98 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Update/word_access_complete/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Update/word_access_complete/word_0/cr
      -- CP-element group 94: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Update/word_access_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_update_start_
      -- 
    cr_2151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(94), ack => array_obj_ref_1122_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1894_elements(98);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	159 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	16 
    -- CP-element group 95: 	33 
    -- CP-element group 95: 	93 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Sample/word_access_start/word_0/$exit
      -- CP-element group 95: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Sample/word_access_start/word_0/ra
      -- CP-element group 95: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Sample/word_access_start/$exit
      -- 
    ra_2141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1122_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (9) 
      -- CP-element group 96: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Update/word_access_complete/word_0/$exit
      -- CP-element group 96: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Update/array_obj_ref_1122_Merge/merge_req
      -- CP-element group 96: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Update/array_obj_ref_1122_Merge/merge_ack
      -- CP-element group 96: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Update/word_access_complete/$exit
      -- CP-element group 96: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Update/word_access_complete/word_0/ca
      -- CP-element group 96: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Update/array_obj_ref_1122_Merge/$entry
      -- CP-element group 96: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_Update/array_obj_ref_1122_Merge/$exit
      -- 
    ca_2152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1122_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	18 
    -- CP-element group 97: 	37 
    -- CP-element group 97: 	96 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_CONTROL_REGISTER_1120_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_CONTROL_REGISTER_1120_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_CONTROL_REGISTER_1120_Sample/req
      -- 
    req_2165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(97), ack => WPIPE_CONTROL_REGISTER_1120_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(18) & SoftwareRegisterAccessDaemon_CP_1894_elements(37) & SoftwareRegisterAccessDaemon_CP_1894_elements(96) & SoftwareRegisterAccessDaemon_CP_1894_elements(99);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	16 
    -- CP-element group 98: 	33 
    -- CP-element group 98: 	94 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_CONTROL_REGISTER_1120_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_CONTROL_REGISTER_1120_update_start_
      -- CP-element group 98: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_CONTROL_REGISTER_1120_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_CONTROL_REGISTER_1120_Sample/ack
      -- CP-element group 98: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_CONTROL_REGISTER_1120_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_CONTROL_REGISTER_1120_Update/req
      -- 
    ack_2166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_CONTROL_REGISTER_1120_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(98)); -- 
    req_2170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(98), ack => WPIPE_CONTROL_REGISTER_1120_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	163 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	97 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_CONTROL_REGISTER_1120_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_CONTROL_REGISTER_1120_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_CONTROL_REGISTER_1120_Update/ack
      -- 
    ack_2171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_CONTROL_REGISTER_1120_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	9 
    -- CP-element group 100: 	18 
    -- CP-element group 100: 	56 
    -- CP-element group 100: marked-predecessors 
    -- CP-element group 100: 	149 
    -- CP-element group 100: 	102 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Sample/word_access_start/$entry
      -- CP-element group 100: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Sample/word_access_start/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Sample/word_access_start/word_0/rr
      -- 
    rr_2188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(100), ack => array_obj_ref_1127_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(9) & SoftwareRegisterAccessDaemon_CP_1894_elements(18) & SoftwareRegisterAccessDaemon_CP_1894_elements(56) & SoftwareRegisterAccessDaemon_CP_1894_elements(149) & SoftwareRegisterAccessDaemon_CP_1894_elements(102);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	110 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_update_start_
      -- CP-element group 101: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Update/$entry
      -- CP-element group 101: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Update/word_access_complete/$entry
      -- CP-element group 101: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Update/word_access_complete/word_0/$entry
      -- CP-element group 101: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Update/word_access_complete/word_0/cr
      -- 
    cr_2199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(101), ack => array_obj_ref_1127_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1894_elements(110);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	160 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	16 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	52 
    -- CP-element group 102:  members (5) 
      -- CP-element group 102: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Sample/word_access_start/$exit
      -- CP-element group 102: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Sample/word_access_start/word_0/$exit
      -- CP-element group 102: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Sample/word_access_start/word_0/ra
      -- 
    ra_2189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1127_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	108 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Update/word_access_complete/$exit
      -- CP-element group 103: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Update/word_access_complete/word_0/$exit
      -- CP-element group 103: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Update/word_access_complete/word_0/ca
      -- CP-element group 103: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Update/array_obj_ref_1127_Merge/$entry
      -- CP-element group 103: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Update/array_obj_ref_1127_Merge/$exit
      -- CP-element group 103: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Update/array_obj_ref_1127_Merge/merge_req
      -- CP-element group 103: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_Update/array_obj_ref_1127_Merge/merge_ack
      -- 
    ca_2200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1127_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	18 
    -- CP-element group 104: 	56 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	106 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1131_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1131_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1131_Sample/req
      -- 
    req_2213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(104), ack => W_update_free_q_pipe_1104_delayed_5_0_1129_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(18) & SoftwareRegisterAccessDaemon_CP_1894_elements(56) & SoftwareRegisterAccessDaemon_CP_1894_elements(106);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	110 
    -- CP-element group 105: 	113 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1131_update_start_
      -- CP-element group 105: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1131_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1131_Update/req
      -- 
    req_2218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(105), ack => W_update_free_q_pipe_1104_delayed_5_0_1129_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(110) & SoftwareRegisterAccessDaemon_CP_1894_elements(113);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106: marked-successors 
    -- CP-element group 106: 	16 
    -- CP-element group 106: 	104 
    -- CP-element group 106: 	52 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1131_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1131_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1131_Sample/ack
      -- 
    ack_2214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_update_free_q_pipe_1104_delayed_5_0_1129_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(106)); -- 
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	112 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1131_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1131_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1131_Update/ack
      -- 
    ack_2219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_update_free_q_pipe_1104_delayed_5_0_1129_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: 	103 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	110 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1138_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1138_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1138_Sample/rr
      -- 
    rr_2227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(108), ack => type_cast_1138_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(107) & SoftwareRegisterAccessDaemon_CP_1894_elements(103) & SoftwareRegisterAccessDaemon_CP_1894_elements(110);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	113 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1138_update_start_
      -- CP-element group 109: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1138_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1138_Update/cr
      -- 
    cr_2232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(109), ack => type_cast_1138_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1894_elements(113);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: 	105 
    -- CP-element group 110: 	101 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1138_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1138_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1138_Sample/ra
      -- 
    ra_2228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1138_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1138_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1138_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/type_cast_1138_Update/ca
      -- 
    ca_2233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1138_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	107 
    -- CP-element group 112: 	111 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	114 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_FREE_Q_1133_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_FREE_Q_1133_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_FREE_Q_1133_Sample/req
      -- 
    req_2241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(112), ack => WPIPE_FREE_Q_1133_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(107) & SoftwareRegisterAccessDaemon_CP_1894_elements(111) & SoftwareRegisterAccessDaemon_CP_1894_elements(114);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113: marked-successors 
    -- CP-element group 113: 	109 
    -- CP-element group 113: 	105 
    -- CP-element group 113:  members (6) 
      -- CP-element group 113: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_FREE_Q_1133_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_FREE_Q_1133_update_start_
      -- CP-element group 113: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_FREE_Q_1133_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_FREE_Q_1133_Sample/ack
      -- CP-element group 113: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_FREE_Q_1133_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_FREE_Q_1133_Update/req
      -- 
    ack_2242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_FREE_Q_1133_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(113)); -- 
    req_2246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(113), ack => WPIPE_FREE_Q_1133_inst_req_1); -- 
    -- CP-element group 114:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	163 
    -- CP-element group 114: marked-successors 
    -- CP-element group 114: 	112 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_FREE_Q_1133_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_FREE_Q_1133_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_FREE_Q_1133_Update/ack
      -- 
    ack_2247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_FREE_Q_1133_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	9 
    -- CP-element group 115: 	18 
    -- CP-element group 115: 	75 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	149 
    -- CP-element group 115: 	117 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Sample/word_access_start/$entry
      -- CP-element group 115: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Sample/word_access_start/word_0/$entry
      -- CP-element group 115: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Sample/word_access_start/word_0/rr
      -- 
    rr_2264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(115), ack => array_obj_ref_1143_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(9) & SoftwareRegisterAccessDaemon_CP_1894_elements(18) & SoftwareRegisterAccessDaemon_CP_1894_elements(75) & SoftwareRegisterAccessDaemon_CP_1894_elements(149) & SoftwareRegisterAccessDaemon_CP_1894_elements(117);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	120 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_update_start_
      -- CP-element group 116: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Update/word_access_complete/$entry
      -- CP-element group 116: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Update/word_access_complete/word_0/$entry
      -- CP-element group 116: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Update/word_access_complete/word_0/cr
      -- 
    cr_2275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(116), ack => array_obj_ref_1143_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1894_elements(120);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	161 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	16 
    -- CP-element group 117: 	115 
    -- CP-element group 117: 	71 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Sample/word_access_start/$exit
      -- CP-element group 117: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Sample/word_access_start/word_0/$exit
      -- CP-element group 117: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Sample/word_access_start/word_0/ra
      -- 
    ra_2265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1143_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (9) 
      -- CP-element group 118: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Update/word_access_complete/$exit
      -- CP-element group 118: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Update/word_access_complete/word_0/$exit
      -- CP-element group 118: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Update/word_access_complete/word_0/ca
      -- CP-element group 118: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Update/array_obj_ref_1143_Merge/$entry
      -- CP-element group 118: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Update/array_obj_ref_1143_Merge/$exit
      -- CP-element group 118: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Update/array_obj_ref_1143_Merge/merge_req
      -- CP-element group 118: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_Update/array_obj_ref_1143_Merge/merge_ack
      -- 
    ca_2276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1143_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	18 
    -- CP-element group 119: 	118 
    -- CP-element group 119: 	75 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	121 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_NUMBER_OF_SERVERS_1141_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_NUMBER_OF_SERVERS_1141_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_NUMBER_OF_SERVERS_1141_Sample/req
      -- 
    req_2289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(119), ack => WPIPE_NUMBER_OF_SERVERS_1141_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 31,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(18) & SoftwareRegisterAccessDaemon_CP_1894_elements(118) & SoftwareRegisterAccessDaemon_CP_1894_elements(75) & SoftwareRegisterAccessDaemon_CP_1894_elements(121);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120: marked-successors 
    -- CP-element group 120: 	16 
    -- CP-element group 120: 	116 
    -- CP-element group 120: 	71 
    -- CP-element group 120:  members (6) 
      -- CP-element group 120: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_NUMBER_OF_SERVERS_1141_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_NUMBER_OF_SERVERS_1141_update_start_
      -- CP-element group 120: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_NUMBER_OF_SERVERS_1141_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_NUMBER_OF_SERVERS_1141_Sample/ack
      -- CP-element group 120: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_NUMBER_OF_SERVERS_1141_Update/$entry
      -- CP-element group 120: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_NUMBER_OF_SERVERS_1141_Update/req
      -- 
    ack_2290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NUMBER_OF_SERVERS_1141_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(120)); -- 
    req_2294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(120), ack => WPIPE_NUMBER_OF_SERVERS_1141_inst_req_1); -- 
    -- CP-element group 121:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	163 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	119 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_NUMBER_OF_SERVERS_1141_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_NUMBER_OF_SERVERS_1141_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_NUMBER_OF_SERVERS_1141_Update/ack
      -- 
    ack_2295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NUMBER_OF_SERVERS_1141_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	9 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	125 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/RPIPE_AFB_NIC_REQUEST_1146_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/RPIPE_AFB_NIC_REQUEST_1146_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/RPIPE_AFB_NIC_REQUEST_1146_Sample/rr
      -- 
    rr_2303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(122), ack => RPIPE_AFB_NIC_REQUEST_1146_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(9) & SoftwareRegisterAccessDaemon_CP_1894_elements(125);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	12 
    -- CP-element group 123: 	124 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	140 
    -- CP-element group 123: 	144 
    -- CP-element group 123: 	132 
    -- CP-element group 123: 	136 
    -- CP-element group 123: 	128 
    -- CP-element group 123: 	152 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/RPIPE_AFB_NIC_REQUEST_1146_update_start_
      -- CP-element group 123: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/RPIPE_AFB_NIC_REQUEST_1146_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/RPIPE_AFB_NIC_REQUEST_1146_Update/cr
      -- 
    cr_2308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(123), ack => RPIPE_AFB_NIC_REQUEST_1146_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(12) & SoftwareRegisterAccessDaemon_CP_1894_elements(124) & SoftwareRegisterAccessDaemon_CP_1894_elements(140) & SoftwareRegisterAccessDaemon_CP_1894_elements(144) & SoftwareRegisterAccessDaemon_CP_1894_elements(132) & SoftwareRegisterAccessDaemon_CP_1894_elements(136) & SoftwareRegisterAccessDaemon_CP_1894_elements(128) & SoftwareRegisterAccessDaemon_CP_1894_elements(152);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	123 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/RPIPE_AFB_NIC_REQUEST_1146_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/RPIPE_AFB_NIC_REQUEST_1146_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/RPIPE_AFB_NIC_REQUEST_1146_Sample/ra
      -- 
    ra_2304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_AFB_NIC_REQUEST_1146_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(124)); -- 
    -- CP-element group 125:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	138 
    -- CP-element group 125: 	142 
    -- CP-element group 125: 	130 
    -- CP-element group 125: 	134 
    -- CP-element group 125: 	150 
    -- CP-element group 125: 	126 
    -- CP-element group 125: marked-successors 
    -- CP-element group 125: 	32 
    -- CP-element group 125: 	122 
    -- CP-element group 125: 	51 
    -- CP-element group 125: 	70 
    -- CP-element group 125:  members (29) 
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/RPIPE_AFB_NIC_REQUEST_1146_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/RPIPE_AFB_NIC_REQUEST_1146_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/RPIPE_AFB_NIC_REQUEST_1146_Update/ca
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_word_address_calculated
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_root_address_calculated
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_offset_calculated
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_index_resized_0
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_index_scaled_0
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_index_computed_0
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_index_resize_0/$entry
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_index_resize_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_index_resize_0/index_resize_req
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_index_resize_0/index_resize_ack
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_index_scale_0/$entry
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_index_scale_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_index_scale_0/scale_rename_req
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_index_scale_0/scale_rename_ack
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_final_index_sum_regn/$entry
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_final_index_sum_regn/$exit
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_final_index_sum_regn/req
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_final_index_sum_regn/ack
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_base_plus_offset/$entry
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_base_plus_offset/$exit
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_base_plus_offset/sum_rename_req
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_base_plus_offset/sum_rename_ack
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_word_addrgen/$entry
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_word_addrgen/$exit
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_word_addrgen/root_register_req
      -- CP-element group 125: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_word_addrgen/root_register_ack
      -- 
    ca_2309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_AFB_NIC_REQUEST_1146_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(125)); -- 
    -- CP-element group 126:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: marked-predecessors 
    -- CP-element group 126: 	128 
    -- CP-element group 126: 	149 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (5) 
      -- CP-element group 126: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Sample/$entry
      -- CP-element group 126: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Sample/word_access_start/$entry
      -- CP-element group 126: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Sample/word_access_start/word_0/$entry
      -- CP-element group 126: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Sample/word_access_start/word_0/rr
      -- 
    rr_2355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(126), ack => array_obj_ref_1199_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(125) & SoftwareRegisterAccessDaemon_CP_1894_elements(128) & SoftwareRegisterAccessDaemon_CP_1894_elements(149);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: marked-predecessors 
    -- CP-element group 127: 	155 
    -- CP-element group 127: 	148 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (5) 
      -- CP-element group 127: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_update_start_
      -- CP-element group 127: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Update/word_access_complete/$entry
      -- CP-element group 127: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Update/word_access_complete/word_0/$entry
      -- CP-element group 127: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Update/word_access_complete/word_0/cr
      -- 
    cr_2366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(127), ack => array_obj_ref_1199_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(155) & SoftwareRegisterAccessDaemon_CP_1894_elements(148);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	162 
    -- CP-element group 128: marked-successors 
    -- CP-element group 128: 	123 
    -- CP-element group 128: 	126 
    -- CP-element group 128:  members (5) 
      -- CP-element group 128: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Sample/word_access_start/$exit
      -- CP-element group 128: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Sample/word_access_start/word_0/$exit
      -- CP-element group 128: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Sample/word_access_start/word_0/ra
      -- 
    ra_2356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1199_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(128)); -- 
    -- CP-element group 129:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	154 
    -- CP-element group 129: 	146 
    -- CP-element group 129:  members (9) 
      -- CP-element group 129: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Update/word_access_complete/$exit
      -- CP-element group 129: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Update/word_access_complete/word_0/$exit
      -- CP-element group 129: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Update/word_access_complete/word_0/ca
      -- CP-element group 129: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Update/array_obj_ref_1199_Merge/$entry
      -- CP-element group 129: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Update/array_obj_ref_1199_Merge/$exit
      -- CP-element group 129: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Update/array_obj_ref_1199_Merge/merge_req
      -- CP-element group 129: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_Update/array_obj_ref_1199_Merge/merge_ack
      -- 
    ca_2367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1199_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(129)); -- 
    -- CP-element group 130:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	125 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	132 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1203_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1203_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1203_Sample/req
      -- 
    req_2380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(130), ack => W_rwbar_1177_delayed_5_0_1201_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(125) & SoftwareRegisterAccessDaemon_CP_1894_elements(132);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	148 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1203_update_start_
      -- CP-element group 131: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1203_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1203_Update/req
      -- 
    req_2385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(131), ack => W_rwbar_1177_delayed_5_0_1201_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1894_elements(148);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: marked-successors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: 	123 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1203_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1203_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1203_Sample/ack
      -- 
    ack_2381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1177_delayed_5_0_1201_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	146 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1203_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1203_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1203_Update/ack
      -- 
    ack_2386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1177_delayed_5_0_1201_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(133)); -- 
    -- CP-element group 134:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	125 
    -- CP-element group 134: marked-predecessors 
    -- CP-element group 134: 	136 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1206_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1206_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1206_Sample/req
      -- 
    req_2394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(134), ack => W_bmask_1178_delayed_5_0_1204_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(125) & SoftwareRegisterAccessDaemon_CP_1894_elements(136);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	148 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1206_update_start_
      -- CP-element group 135: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1206_Update/$entry
      -- CP-element group 135: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1206_Update/req
      -- 
    req_2399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(135), ack => W_bmask_1178_delayed_5_0_1204_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1894_elements(148);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: marked-successors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: 	123 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1206_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1206_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1206_Sample/ack
      -- 
    ack_2395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_1178_delayed_5_0_1204_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	146 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1206_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1206_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1206_Update/ack
      -- 
    ack_2400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_1178_delayed_5_0_1204_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(137)); -- 
    -- CP-element group 138:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	125 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	140 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1209_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1209_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1209_Sample/req
      -- 
    req_2408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(138), ack => W_wdata_1180_delayed_5_0_1207_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(125) & SoftwareRegisterAccessDaemon_CP_1894_elements(140);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	148 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1209_update_start_
      -- CP-element group 139: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1209_Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1209_Update/req
      -- 
    req_2413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(139), ack => W_wdata_1180_delayed_5_0_1207_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1894_elements(148);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140: marked-successors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: 	123 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1209_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1209_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1209_Sample/ack
      -- 
    ack_2409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_1180_delayed_5_0_1207_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	146 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1209_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1209_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1209_Update/ack
      -- 
    ack_2414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_1180_delayed_5_0_1207_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(141)); -- 
    -- CP-element group 142:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	125 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	144 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1212_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1212_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1212_Sample/req
      -- 
    req_2422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(142), ack => W_index_1181_delayed_5_0_1210_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(125) & SoftwareRegisterAccessDaemon_CP_1894_elements(144);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	148 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1212_update_start_
      -- CP-element group 143: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1212_Update/$entry
      -- CP-element group 143: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1212_Update/req
      -- 
    req_2427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(143), ack => W_index_1181_delayed_5_0_1210_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1894_elements(148);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: marked-successors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: 	123 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1212_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1212_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1212_Sample/ack
      -- 
    ack_2423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_1181_delayed_5_0_1210_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1212_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1212_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1212_Update/ack
      -- 
    ack_2428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_1181_delayed_5_0_1210_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(145)); -- 
    -- CP-element group 146:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	141 
    -- CP-element group 146: 	145 
    -- CP-element group 146: 	133 
    -- CP-element group 146: 	137 
    -- CP-element group 146: 	158 
    -- CP-element group 146: 	159 
    -- CP-element group 146: 	160 
    -- CP-element group 146: 	161 
    -- CP-element group 146: 	162 
    -- CP-element group 146: 	129 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	148 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/call_stmt_1219_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/call_stmt_1219_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/call_stmt_1219_Sample/crr
      -- 
    crr_2436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(146), ack => call_stmt_1219_call_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 31,5 => 31,6 => 31,7 => 31,8 => 31,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 1);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(141) & SoftwareRegisterAccessDaemon_CP_1894_elements(145) & SoftwareRegisterAccessDaemon_CP_1894_elements(133) & SoftwareRegisterAccessDaemon_CP_1894_elements(137) & SoftwareRegisterAccessDaemon_CP_1894_elements(158) & SoftwareRegisterAccessDaemon_CP_1894_elements(159) & SoftwareRegisterAccessDaemon_CP_1894_elements(160) & SoftwareRegisterAccessDaemon_CP_1894_elements(161) & SoftwareRegisterAccessDaemon_CP_1894_elements(162) & SoftwareRegisterAccessDaemon_CP_1894_elements(129) & SoftwareRegisterAccessDaemon_CP_1894_elements(148);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	149 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/call_stmt_1219_update_start_
      -- CP-element group 147: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/call_stmt_1219_Update/$entry
      -- CP-element group 147: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/call_stmt_1219_Update/ccr
      -- 
    ccr_2441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(147), ack => call_stmt_1219_call_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1894_elements(149);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	139 
    -- CP-element group 148: 	143 
    -- CP-element group 148: 	131 
    -- CP-element group 148: 	135 
    -- CP-element group 148: 	146 
    -- CP-element group 148: 	127 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/call_stmt_1219_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/call_stmt_1219_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/call_stmt_1219_Sample/cra
      -- 
    cra_2437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1219_call_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(148)); -- 
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	163 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: 	115 
    -- CP-element group 149: 	126 
    -- CP-element group 149: 	93 
    -- CP-element group 149: 	100 
    -- CP-element group 149: 	89 
    -- CP-element group 149:  members (4) 
      -- CP-element group 149: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/call_stmt_1219_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/call_stmt_1219_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/call_stmt_1219_Update/cca
      -- CP-element group 149: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/ring_reenable_memory_space_0
      -- 
    cca_2442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1219_call_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(149)); -- 
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	125 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1222_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1222_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1222_Sample/req
      -- 
    req_2450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(150), ack => W_rwbar_1185_delayed_5_0_1220_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(125) & SoftwareRegisterAccessDaemon_CP_1894_elements(152);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	155 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1222_update_start_
      -- CP-element group 151: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1222_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1222_Update/req
      -- 
    req_2455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(151), ack => W_rwbar_1185_delayed_5_0_1220_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1894_elements(155);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	123 
    -- CP-element group 152: 	150 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1222_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1222_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1222_Sample/ack
      -- 
    ack_2451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1185_delayed_5_0_1220_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1222_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1222_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/assign_stmt_1222_Update/ack
      -- 
    ack_2456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1185_delayed_5_0_1220_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	129 
    -- CP-element group 154: 	153 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_AFB_NIC_RESPONSE_1236_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_AFB_NIC_RESPONSE_1236_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_AFB_NIC_RESPONSE_1236_Sample/req
      -- 
    req_2464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(154), ack => WPIPE_AFB_NIC_RESPONSE_1236_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(129) & SoftwareRegisterAccessDaemon_CP_1894_elements(153) & SoftwareRegisterAccessDaemon_CP_1894_elements(156);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	151 
    -- CP-element group 155: 	127 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_AFB_NIC_RESPONSE_1236_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_AFB_NIC_RESPONSE_1236_update_start_
      -- CP-element group 155: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_AFB_NIC_RESPONSE_1236_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_AFB_NIC_RESPONSE_1236_Sample/ack
      -- CP-element group 155: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_AFB_NIC_RESPONSE_1236_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_AFB_NIC_RESPONSE_1236_Update/req
      -- 
    ack_2465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_AFB_NIC_RESPONSE_1236_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(155)); -- 
    req_2469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1894_elements(155), ack => WPIPE_AFB_NIC_RESPONSE_1236_inst_req_1); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	163 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_AFB_NIC_RESPONSE_1236_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_AFB_NIC_RESPONSE_1236_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/WPIPE_AFB_NIC_RESPONSE_1236_Update/ack
      -- 
    ack_2470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_AFB_NIC_RESPONSE_1236_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(156)); -- 
    -- CP-element group 157:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	9 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	10 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(157) is a control-delay.
    cp_element_157_delay: control_delay_element  generic map(name => " 157_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1894_elements(9), ack => SoftwareRegisterAccessDaemon_CP_1894_elements(157), clk => clk, reset =>reset);
    -- CP-element group 158:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	91 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	146 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1091_call_stmt_1219_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(158) is a control-delay.
    cp_element_158_delay: control_delay_element  generic map(name => " 158_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1894_elements(91), ack => SoftwareRegisterAccessDaemon_CP_1894_elements(158), clk => clk, reset =>reset);
    -- CP-element group 159:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	95 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	146 
    -- CP-element group 159:  members (1) 
      -- CP-element group 159: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1122_call_stmt_1219_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(159) is a control-delay.
    cp_element_159_delay: control_delay_element  generic map(name => " 159_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1894_elements(95), ack => SoftwareRegisterAccessDaemon_CP_1894_elements(159), clk => clk, reset =>reset);
    -- CP-element group 160:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	102 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	146 
    -- CP-element group 160:  members (1) 
      -- CP-element group 160: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1127_call_stmt_1219_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(160) is a control-delay.
    cp_element_160_delay: control_delay_element  generic map(name => " 160_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1894_elements(102), ack => SoftwareRegisterAccessDaemon_CP_1894_elements(160), clk => clk, reset =>reset);
    -- CP-element group 161:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	117 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	146 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1143_call_stmt_1219_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(161) is a control-delay.
    cp_element_161_delay: control_delay_element  generic map(name => " 161_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1894_elements(117), ack => SoftwareRegisterAccessDaemon_CP_1894_elements(161), clk => clk, reset =>reset);
    -- CP-element group 162:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	128 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	146 
    -- CP-element group 162:  members (1) 
      -- CP-element group 162: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/array_obj_ref_1199_call_stmt_1219_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1894_elements(162) is a control-delay.
    cp_element_162_delay: control_delay_element  generic map(name => " 162_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1894_elements(128), ack => SoftwareRegisterAccessDaemon_CP_1894_elements(162), clk => clk, reset =>reset);
    -- CP-element group 163:  join  transition  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	12 
    -- CP-element group 163: 	121 
    -- CP-element group 163: 	156 
    -- CP-element group 163: 	149 
    -- CP-element group 163: 	92 
    -- CP-element group 163: 	114 
    -- CP-element group 163: 	99 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	6 
    -- CP-element group 163:  members (1) 
      -- CP-element group 163: 	 branch_block_stmt_1063/do_while_stmt_1064/do_while_stmt_1064_loop_body/$exit
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 31,1 => 31,2 => 31,3 => 31,4 => 31,5 => 31,6 => 31);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1894_elements(12) & SoftwareRegisterAccessDaemon_CP_1894_elements(121) & SoftwareRegisterAccessDaemon_CP_1894_elements(156) & SoftwareRegisterAccessDaemon_CP_1894_elements(149) & SoftwareRegisterAccessDaemon_CP_1894_elements(92) & SoftwareRegisterAccessDaemon_CP_1894_elements(114) & SoftwareRegisterAccessDaemon_CP_1894_elements(99);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	5 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_1063/do_while_stmt_1064/loop_exit/$exit
      -- CP-element group 164: 	 branch_block_stmt_1063/do_while_stmt_1064/loop_exit/ack
      -- 
    ack_2481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1064_branch_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	5 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (2) 
      -- CP-element group 165: 	 branch_block_stmt_1063/do_while_stmt_1064/loop_taken/$exit
      -- CP-element group 165: 	 branch_block_stmt_1063/do_while_stmt_1064/loop_taken/ack
      -- 
    ack_2485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1064_branch_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1894_elements(165)); -- 
    -- CP-element group 166:  transition  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	3 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	1 
    -- CP-element group 166:  members (1) 
      -- CP-element group 166: 	 branch_block_stmt_1063/do_while_stmt_1064/$exit
      -- 
    SoftwareRegisterAccessDaemon_CP_1894_elements(166) <= SoftwareRegisterAccessDaemon_CP_1894_elements(3);
    SoftwareRegisterAccessDaemon_do_while_stmt_1064_terminator_2486: loop_terminator -- 
      generic map (name => " SoftwareRegisterAccessDaemon_do_while_stmt_1064_terminator_2486", max_iterations_in_flight =>31) 
      port map(loop_body_exit => SoftwareRegisterAccessDaemon_CP_1894_elements(6),loop_continue => SoftwareRegisterAccessDaemon_CP_1894_elements(165),loop_terminate => SoftwareRegisterAccessDaemon_CP_1894_elements(164),loop_back => SoftwareRegisterAccessDaemon_CP_1894_elements(4),loop_exit => SoftwareRegisterAccessDaemon_CP_1894_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1066_phi_seq_1957_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(21);
      SoftwareRegisterAccessDaemon_CP_1894_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(24);
      SoftwareRegisterAccessDaemon_CP_1894_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(26);
      SoftwareRegisterAccessDaemon_CP_1894_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(19);
      SoftwareRegisterAccessDaemon_CP_1894_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(28);
      SoftwareRegisterAccessDaemon_CP_1894_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(30);
      SoftwareRegisterAccessDaemon_CP_1894_elements(20) <= phi_mux_reqs(1);
      phi_stmt_1066_phi_seq_1957 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1066_phi_seq_1957") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_1894_elements(11), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_1894_elements(17), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_1894_elements(13), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_1894_elements(18), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_1894_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1072_phi_seq_2001_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(40);
      SoftwareRegisterAccessDaemon_CP_1894_elements(43)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(43);
      SoftwareRegisterAccessDaemon_CP_1894_elements(44)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(45);
      SoftwareRegisterAccessDaemon_CP_1894_elements(41) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(38);
      SoftwareRegisterAccessDaemon_CP_1894_elements(47)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(49);
      SoftwareRegisterAccessDaemon_CP_1894_elements(48)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(50);
      SoftwareRegisterAccessDaemon_CP_1894_elements(39) <= phi_mux_reqs(1);
      phi_stmt_1072_phi_seq_2001 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1072_phi_seq_2001") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_1894_elements(34), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_1894_elements(35), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_1894_elements(36), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_1894_elements(37), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_1894_elements(42), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1077_phi_seq_2045_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(59);
      SoftwareRegisterAccessDaemon_CP_1894_elements(62)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(62);
      SoftwareRegisterAccessDaemon_CP_1894_elements(63)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(64);
      SoftwareRegisterAccessDaemon_CP_1894_elements(60) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(57);
      SoftwareRegisterAccessDaemon_CP_1894_elements(66)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(68);
      SoftwareRegisterAccessDaemon_CP_1894_elements(67)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(69);
      SoftwareRegisterAccessDaemon_CP_1894_elements(58) <= phi_mux_reqs(1);
      phi_stmt_1077_phi_seq_2045 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1077_phi_seq_2045") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_1894_elements(53), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_1894_elements(54), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_1894_elements(55), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_1894_elements(56), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_1894_elements(61), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1082_phi_seq_2089_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(78);
      SoftwareRegisterAccessDaemon_CP_1894_elements(81)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(81);
      SoftwareRegisterAccessDaemon_CP_1894_elements(82)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(83);
      SoftwareRegisterAccessDaemon_CP_1894_elements(79) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(76);
      SoftwareRegisterAccessDaemon_CP_1894_elements(85)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(87);
      SoftwareRegisterAccessDaemon_CP_1894_elements(86)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(88);
      SoftwareRegisterAccessDaemon_CP_1894_elements(77) <= phi_mux_reqs(1);
      phi_stmt_1082_phi_seq_2089 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1082_phi_seq_2089") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_1894_elements(72), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_1894_elements(73), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_1894_elements(74), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_1894_elements(75), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_1894_elements(80), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1919_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(7);
        preds(1)  <= SoftwareRegisterAccessDaemon_CP_1894_elements(8);
        entry_tmerge_1919 : transition_merge -- 
          generic map(name => " entry_tmerge_1919")
          port map (preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1894_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_1100_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1108_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1116_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u32_u35_1137_wire : std_logic_vector(34 downto 0);
    signal EQ_u1_u1_1176_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_1185_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_1194_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_1173_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_1182_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_1191_wire : std_logic_vector(0 downto 0);
    signal FREE_Q_32_1128 : std_logic_vector(31 downto 0);
    signal INIT_1066 : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1097_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1105_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1113_wire : std_logic_vector(0 downto 0);
    signal R_index_1198_resized : std_logic_vector(5 downto 0);
    signal R_index_1198_scaled : std_logic_vector(5 downto 0);
    signal addr_1161 : std_logic_vector(35 downto 0);
    signal array_obj_ref_1091_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1091_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1122_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1122_wire : std_logic_vector(31 downto 0);
    signal array_obj_ref_1122_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1127_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1127_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1143_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1143_wire : std_logic_vector(31 downto 0);
    signal array_obj_ref_1143_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1199_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1199_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_1199_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1199_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_1199_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_1199_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1199_word_offset_0 : std_logic_vector(5 downto 0);
    signal bmask_1157 : std_logic_vector(3 downto 0);
    signal bmask_1178_delayed_5_0_1206 : std_logic_vector(3 downto 0);
    signal check_control_regsiter_1178 : std_logic_vector(0 downto 0);
    signal check_control_regsiter_1178_1076_buffered : std_logic_vector(0 downto 0);
    signal check_free_q_1187 : std_logic_vector(0 downto 0);
    signal check_free_q_1187_1081_buffered : std_logic_vector(0 downto 0);
    signal check_num_server_1196 : std_logic_vector(0 downto 0);
    signal check_num_server_1196_1086_buffered : std_logic_vector(0 downto 0);
    signal control_data_1092 : std_logic_vector(31 downto 0);
    signal control_register_1072 : std_logic_vector(0 downto 0);
    signal free_q_1077 : std_logic_vector(0 downto 0);
    signal index_1169 : std_logic_vector(5 downto 0);
    signal index_1181_delayed_5_0_1212 : std_logic_vector(5 downto 0);
    signal konst_1172_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1175_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1181_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1184_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1190_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1193_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1240_wire_constant : std_logic_vector(0 downto 0);
    signal num_server_1082 : std_logic_vector(0 downto 0);
    signal rdata_1229 : std_logic_vector(31 downto 0);
    signal req_1147 : std_logic_vector(73 downto 0);
    signal resp_1235 : std_logic_vector(32 downto 0);
    signal rval_1200 : std_logic_vector(31 downto 0);
    signal rwbar_1153 : std_logic_vector(0 downto 0);
    signal rwbar_1177_delayed_5_0_1203 : std_logic_vector(0 downto 0);
    signal rwbar_1185_delayed_5_0_1222 : std_logic_vector(0 downto 0);
    signal type_cast_1069_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1071_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1075_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1080_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1085_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1136_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_1138_wire : std_logic_vector(35 downto 0);
    signal type_cast_1227_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1232_wire_constant : std_logic_vector(0 downto 0);
    signal update_control_register_pipe_1102 : std_logic_vector(0 downto 0);
    signal update_free_q_pipe_1104_delayed_5_0_1131 : std_logic_vector(0 downto 0);
    signal update_free_q_pipe_1110 : std_logic_vector(0 downto 0);
    signal update_server_num_1118 : std_logic_vector(0 downto 0);
    signal wdata_1165 : std_logic_vector(31 downto 0);
    signal wdata_1180_delayed_5_0_1209 : std_logic_vector(31 downto 0);
    signal wval_1219 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1091_word_address_0 <= "000000";
    array_obj_ref_1122_word_address_0 <= "000000";
    array_obj_ref_1127_word_address_0 <= "010010";
    array_obj_ref_1143_word_address_0 <= "000001";
    array_obj_ref_1199_offset_scale_factor_0 <= "000001";
    array_obj_ref_1199_resized_base_address <= "000000";
    array_obj_ref_1199_word_offset_0 <= "000000";
    konst_1172_wire_constant <= "000000";
    konst_1175_wire_constant <= "0";
    konst_1181_wire_constant <= "010010";
    konst_1184_wire_constant <= "0";
    konst_1190_wire_constant <= "000001";
    konst_1193_wire_constant <= "0";
    konst_1240_wire_constant <= "1";
    type_cast_1069_wire_constant <= "0";
    type_cast_1071_wire_constant <= "1";
    type_cast_1075_wire_constant <= "0";
    type_cast_1080_wire_constant <= "0";
    type_cast_1085_wire_constant <= "0";
    type_cast_1136_wire_constant <= "000";
    type_cast_1227_wire_constant <= "00000000000000000000000000000000";
    type_cast_1232_wire_constant <= "0";
    phi_stmt_1066: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1069_wire_constant & type_cast_1071_wire_constant;
      req <= phi_stmt_1066_req_0 & phi_stmt_1066_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1066",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1066_ack_0,
          idata => idata,
          odata => INIT_1066,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1066
    phi_stmt_1072: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1075_wire_constant & check_control_regsiter_1178_1076_buffered;
      req <= phi_stmt_1072_req_0 & phi_stmt_1072_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1072",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1072_ack_0,
          idata => idata,
          odata => control_register_1072,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1072
    phi_stmt_1077: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1080_wire_constant & check_free_q_1187_1081_buffered;
      req <= phi_stmt_1077_req_0 & phi_stmt_1077_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1077",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1077_ack_0,
          idata => idata,
          odata => free_q_1077,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1077
    phi_stmt_1082: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1085_wire_constant & check_num_server_1196_1086_buffered;
      req <= phi_stmt_1082_req_0 & phi_stmt_1082_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1082",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1082_ack_0,
          idata => idata,
          odata => num_server_1082,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1082
    -- flow-through select operator MUX_1228_inst
    rdata_1229 <= rval_1200 when (rwbar_1185_delayed_5_0_1222(0) /=  '0') else type_cast_1227_wire_constant;
    -- flow-through slice operator slice_1152_inst
    rwbar_1153 <= req_1147(72 downto 72);
    -- flow-through slice operator slice_1156_inst
    bmask_1157 <= req_1147(71 downto 68);
    -- flow-through slice operator slice_1160_inst
    addr_1161 <= req_1147(67 downto 32);
    -- flow-through slice operator slice_1164_inst
    wdata_1165 <= req_1147(31 downto 0);
    -- flow-through slice operator slice_1168_inst
    index_1169 <= addr_1161(7 downto 2);
    W_bmask_1178_delayed_5_0_1204_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_bmask_1178_delayed_5_0_1204_inst_req_0;
      W_bmask_1178_delayed_5_0_1204_inst_ack_0<= wack(0);
      rreq(0) <= W_bmask_1178_delayed_5_0_1204_inst_req_1;
      W_bmask_1178_delayed_5_0_1204_inst_ack_1<= rack(0);
      W_bmask_1178_delayed_5_0_1204_inst : InterlockBuffer generic map ( -- 
        name => "W_bmask_1178_delayed_5_0_1204_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => bmask_1157,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => bmask_1178_delayed_5_0_1206,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_index_1181_delayed_5_0_1210_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_index_1181_delayed_5_0_1210_inst_req_0;
      W_index_1181_delayed_5_0_1210_inst_ack_0<= wack(0);
      rreq(0) <= W_index_1181_delayed_5_0_1210_inst_req_1;
      W_index_1181_delayed_5_0_1210_inst_ack_1<= rack(0);
      W_index_1181_delayed_5_0_1210_inst : InterlockBuffer generic map ( -- 
        name => "W_index_1181_delayed_5_0_1210_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => index_1169,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => index_1181_delayed_5_0_1212,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_1177_delayed_5_0_1201_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_1177_delayed_5_0_1201_inst_req_0;
      W_rwbar_1177_delayed_5_0_1201_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_1177_delayed_5_0_1201_inst_req_1;
      W_rwbar_1177_delayed_5_0_1201_inst_ack_1<= rack(0);
      W_rwbar_1177_delayed_5_0_1201_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_1177_delayed_5_0_1201_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_1153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_1177_delayed_5_0_1203,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_1185_delayed_5_0_1220_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_1185_delayed_5_0_1220_inst_req_0;
      W_rwbar_1185_delayed_5_0_1220_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_1185_delayed_5_0_1220_inst_req_1;
      W_rwbar_1185_delayed_5_0_1220_inst_ack_1<= rack(0);
      W_rwbar_1185_delayed_5_0_1220_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_1185_delayed_5_0_1220_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_1153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_1185_delayed_5_0_1222,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_update_free_q_pipe_1104_delayed_5_0_1129_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_update_free_q_pipe_1104_delayed_5_0_1129_inst_req_0;
      W_update_free_q_pipe_1104_delayed_5_0_1129_inst_ack_0<= wack(0);
      rreq(0) <= W_update_free_q_pipe_1104_delayed_5_0_1129_inst_req_1;
      W_update_free_q_pipe_1104_delayed_5_0_1129_inst_ack_1<= rack(0);
      W_update_free_q_pipe_1104_delayed_5_0_1129_inst : InterlockBuffer generic map ( -- 
        name => "W_update_free_q_pipe_1104_delayed_5_0_1129_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => update_free_q_pipe_1110,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => update_free_q_pipe_1104_delayed_5_0_1131,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_wdata_1180_delayed_5_0_1207_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_wdata_1180_delayed_5_0_1207_inst_req_0;
      W_wdata_1180_delayed_5_0_1207_inst_ack_0<= wack(0);
      rreq(0) <= W_wdata_1180_delayed_5_0_1207_inst_req_1;
      W_wdata_1180_delayed_5_0_1207_inst_ack_1<= rack(0);
      W_wdata_1180_delayed_5_0_1207_inst : InterlockBuffer generic map ( -- 
        name => "W_wdata_1180_delayed_5_0_1207_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => wdata_1165,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => wdata_1180_delayed_5_0_1209,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    check_control_regsiter_1178_1076_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= check_control_regsiter_1178_1076_buf_req_0;
      check_control_regsiter_1178_1076_buf_ack_0<= wack(0);
      rreq(0) <= check_control_regsiter_1178_1076_buf_req_1;
      check_control_regsiter_1178_1076_buf_ack_1<= rack(0);
      check_control_regsiter_1178_1076_buf : InterlockBuffer generic map ( -- 
        name => "check_control_regsiter_1178_1076_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => check_control_regsiter_1178,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => check_control_regsiter_1178_1076_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    check_free_q_1187_1081_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= check_free_q_1187_1081_buf_req_0;
      check_free_q_1187_1081_buf_ack_0<= wack(0);
      rreq(0) <= check_free_q_1187_1081_buf_req_1;
      check_free_q_1187_1081_buf_ack_1<= rack(0);
      check_free_q_1187_1081_buf : InterlockBuffer generic map ( -- 
        name => "check_free_q_1187_1081_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => check_free_q_1187,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => check_free_q_1187_1081_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    check_num_server_1196_1086_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= check_num_server_1196_1086_buf_req_0;
      check_num_server_1196_1086_buf_ack_0<= wack(0);
      rreq(0) <= check_num_server_1196_1086_buf_req_1;
      check_num_server_1196_1086_buf_ack_1<= rack(0);
      check_num_server_1196_1086_buf : InterlockBuffer generic map ( -- 
        name => "check_num_server_1196_1086_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => check_num_server_1196,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => check_num_server_1196_1086_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1138_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1138_inst_req_0;
      type_cast_1138_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1138_inst_req_1;
      type_cast_1138_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  update_free_q_pipe_1104_delayed_5_0_1131(0);
      type_cast_1138_inst_gI: SplitGuardInterface generic map(name => "type_cast_1138_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1138_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1138_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 35,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => CONCAT_u32_u35_1137_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1138_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1091_gather_scatter
    process(array_obj_ref_1091_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1091_data_0;
      ov(31 downto 0) := iv;
      control_data_1092 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1122_gather_scatter
    process(array_obj_ref_1122_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1122_data_0;
      ov(31 downto 0) := iv;
      array_obj_ref_1122_wire <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1127_gather_scatter
    process(array_obj_ref_1127_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1127_data_0;
      ov(31 downto 0) := iv;
      FREE_Q_32_1128 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1143_gather_scatter
    process(array_obj_ref_1143_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1143_data_0;
      ov(31 downto 0) := iv;
      array_obj_ref_1143_wire <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1199_addr_0
    process(array_obj_ref_1199_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1199_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_1199_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1199_gather_scatter
    process(array_obj_ref_1199_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1199_data_0;
      ov(31 downto 0) := iv;
      rval_1200 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1199_index_0_rename
    process(R_index_1198_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_1198_resized;
      ov(5 downto 0) := iv;
      R_index_1198_scaled <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1199_index_0_resize
    process(index_1169) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_1169;
      ov(5 downto 0) := iv;
      R_index_1198_resized <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1199_index_offset
    process(R_index_1198_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_1198_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_1199_final_offset <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1199_root_address_inst
    process(array_obj_ref_1199_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1199_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_1199_root_address <= ov(5 downto 0);
      --
    end process;
    do_while_stmt_1064_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1240_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1064_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1064_branch_req_0,
          ack0 => do_while_stmt_1064_branch_ack_0,
          ack1 => do_while_stmt_1064_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_1100_inst
    process(INIT_1066, control_register_1072) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(INIT_1066, control_register_1072, tmp_var);
      AND_u1_u1_1100_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1108_inst
    process(INIT_1066, free_q_1077) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(INIT_1066, free_q_1077, tmp_var);
      AND_u1_u1_1108_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1116_inst
    process(INIT_1066, num_server_1082) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(INIT_1066, num_server_1082, tmp_var);
      AND_u1_u1_1116_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1177_inst
    process(EQ_u6_u1_1173_wire, EQ_u1_u1_1176_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u6_u1_1173_wire, EQ_u1_u1_1176_wire, tmp_var);
      check_control_regsiter_1178 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1186_inst
    process(EQ_u6_u1_1182_wire, EQ_u1_u1_1185_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u6_u1_1182_wire, EQ_u1_u1_1185_wire, tmp_var);
      check_free_q_1187 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1195_inst
    process(EQ_u6_u1_1191_wire, EQ_u1_u1_1194_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u6_u1_1191_wire, EQ_u1_u1_1194_wire, tmp_var);
      check_num_server_1196 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u33_1234_inst
    process(type_cast_1232_wire_constant, rdata_1229) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1232_wire_constant, rdata_1229, tmp_var);
      resp_1235 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u35_1137_inst
    process(FREE_Q_32_1128) -- 
      variable tmp_var : std_logic_vector(34 downto 0); -- 
    begin -- 
      ApConcat_proc(FREE_Q_32_1128, type_cast_1136_wire_constant, tmp_var);
      CONCAT_u32_u35_1137_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1176_inst
    process(rwbar_1153) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rwbar_1153, konst_1175_wire_constant, tmp_var);
      EQ_u1_u1_1176_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1185_inst
    process(rwbar_1153) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rwbar_1153, konst_1184_wire_constant, tmp_var);
      EQ_u1_u1_1185_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1194_inst
    process(rwbar_1153) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rwbar_1153, konst_1193_wire_constant, tmp_var);
      EQ_u1_u1_1194_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u6_u1_1173_inst
    process(index_1169) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_1169, konst_1172_wire_constant, tmp_var);
      EQ_u6_u1_1173_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u6_u1_1182_inst
    process(index_1169) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_1169, konst_1181_wire_constant, tmp_var);
      EQ_u6_u1_1182_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u6_u1_1191_inst
    process(index_1169) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_1169, konst_1190_wire_constant, tmp_var);
      EQ_u6_u1_1191_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1097_inst
    process(INIT_1066) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", INIT_1066, tmp_var);
      NOT_u1_u1_1097_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1105_inst
    process(INIT_1066) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", INIT_1066, tmp_var);
      NOT_u1_u1_1105_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1113_inst
    process(INIT_1066) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", INIT_1066, tmp_var);
      NOT_u1_u1_1113_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1101_inst
    process(NOT_u1_u1_1097_wire, AND_u1_u1_1100_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1097_wire, AND_u1_u1_1100_wire, tmp_var);
      update_control_register_pipe_1102 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1109_inst
    process(NOT_u1_u1_1105_wire, AND_u1_u1_1108_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1105_wire, AND_u1_u1_1108_wire, tmp_var);
      update_free_q_pipe_1110 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1117_inst
    process(NOT_u1_u1_1113_wire, AND_u1_u1_1116_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1113_wire, AND_u1_u1_1116_wire, tmp_var);
      update_server_num_1118 <= tmp_var; --
    end process;
    -- shared load operator group (0) : array_obj_ref_1199_load_0 array_obj_ref_1143_load_0 array_obj_ref_1127_load_0 array_obj_ref_1122_load_0 array_obj_ref_1091_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(29 downto 0);
      signal data_out: std_logic_vector(159 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 4 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 4 downto 0);
      signal guard_vector : std_logic_vector( 4 downto 0);
      constant inBUFs : IntegerArray(4 downto 0) := (4 => 2, 3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(4 downto 0) := (4 => 2, 3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(4 downto 0) := (0 => false, 1 => true, 2 => true, 3 => true, 4 => false);
      constant guardBuffering: IntegerArray(4 downto 0)  := (0 => 5, 1 => 5, 2 => 5, 3 => 5, 4 => 5);
      -- 
    begin -- 
      reqL_unguarded(4) <= array_obj_ref_1199_load_0_req_0;
      reqL_unguarded(3) <= array_obj_ref_1143_load_0_req_0;
      reqL_unguarded(2) <= array_obj_ref_1127_load_0_req_0;
      reqL_unguarded(1) <= array_obj_ref_1122_load_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_1091_load_0_req_0;
      array_obj_ref_1199_load_0_ack_0 <= ackL_unguarded(4);
      array_obj_ref_1143_load_0_ack_0 <= ackL_unguarded(3);
      array_obj_ref_1127_load_0_ack_0 <= ackL_unguarded(2);
      array_obj_ref_1122_load_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_1091_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(4) <= array_obj_ref_1199_load_0_req_1;
      reqR_unguarded(3) <= array_obj_ref_1143_load_0_req_1;
      reqR_unguarded(2) <= array_obj_ref_1127_load_0_req_1;
      reqR_unguarded(1) <= array_obj_ref_1122_load_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_1091_load_0_req_1;
      array_obj_ref_1199_load_0_ack_1 <= ackR_unguarded(4);
      array_obj_ref_1143_load_0_ack_1 <= ackR_unguarded(3);
      array_obj_ref_1127_load_0_ack_1 <= ackR_unguarded(2);
      array_obj_ref_1122_load_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_1091_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <= update_control_register_pipe_1102(0);
      guard_vector(2)  <= update_free_q_pipe_1110(0);
      guard_vector(3)  <= update_server_num_1118(0);
      guard_vector(4)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 5, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_1199_word_address_0 & array_obj_ref_1143_word_address_0 & array_obj_ref_1127_word_address_0 & array_obj_ref_1122_word_address_0 & array_obj_ref_1091_word_address_0;
      array_obj_ref_1199_data_0 <= data_out(159 downto 128);
      array_obj_ref_1143_data_0 <= data_out(127 downto 96);
      array_obj_ref_1127_data_0 <= data_out(95 downto 64);
      array_obj_ref_1122_data_0 <= data_out(63 downto 32);
      array_obj_ref_1091_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 6,
        num_reqs => 5,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(5 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 5,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_AFB_NIC_REQUEST_1146_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(73 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_AFB_NIC_REQUEST_1146_inst_req_0;
      RPIPE_AFB_NIC_REQUEST_1146_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_AFB_NIC_REQUEST_1146_inst_req_1;
      RPIPE_AFB_NIC_REQUEST_1146_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      req_1147 <= data_out(73 downto 0);
      AFB_NIC_REQUEST_read_0_gI: SplitGuardInterface generic map(name => "AFB_NIC_REQUEST_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      AFB_NIC_REQUEST_read_0: InputPortRevised -- 
        generic map ( name => "AFB_NIC_REQUEST_read_0", data_width => 74,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => AFB_NIC_REQUEST_pipe_read_req(0),
          oack => AFB_NIC_REQUEST_pipe_read_ack(0),
          odata => AFB_NIC_REQUEST_pipe_read_data(73 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_AFB_NIC_RESPONSE_1236_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_AFB_NIC_RESPONSE_1236_inst_req_0;
      WPIPE_AFB_NIC_RESPONSE_1236_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_AFB_NIC_RESPONSE_1236_inst_req_1;
      WPIPE_AFB_NIC_RESPONSE_1236_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= resp_1235;
      AFB_NIC_RESPONSE_write_0_gI: SplitGuardInterface generic map(name => "AFB_NIC_RESPONSE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      AFB_NIC_RESPONSE_write_0: OutputPortRevised -- 
        generic map ( name => "AFB_NIC_RESPONSE", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => AFB_NIC_RESPONSE_pipe_write_req(0),
          oack => AFB_NIC_RESPONSE_pipe_write_ack(0),
          odata => AFB_NIC_RESPONSE_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_CONTROL_REGISTER_1120_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_CONTROL_REGISTER_1120_inst_req_0;
      WPIPE_CONTROL_REGISTER_1120_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_CONTROL_REGISTER_1120_inst_req_1;
      WPIPE_CONTROL_REGISTER_1120_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_control_register_pipe_1102(0);
      data_in <= array_obj_ref_1122_wire;
      CONTROL_REGISTER_write_1_gI: SplitGuardInterface generic map(name => "CONTROL_REGISTER_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      CONTROL_REGISTER_write_1: OutputPortRevised -- 
        generic map ( name => "CONTROL_REGISTER", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => CONTROL_REGISTER_pipe_write_req(0),
          oack => CONTROL_REGISTER_pipe_write_ack(0),
          odata => CONTROL_REGISTER_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_FREE_Q_1133_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_FREE_Q_1133_inst_req_0;
      WPIPE_FREE_Q_1133_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_FREE_Q_1133_inst_req_1;
      WPIPE_FREE_Q_1133_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_free_q_pipe_1104_delayed_5_0_1131(0);
      data_in <= type_cast_1138_wire;
      FREE_Q_write_2_gI: SplitGuardInterface generic map(name => "FREE_Q_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      FREE_Q_write_2: OutputPortRevised -- 
        generic map ( name => "FREE_Q", data_width => 36, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => FREE_Q_pipe_write_req(0),
          oack => FREE_Q_pipe_write_ack(0),
          odata => FREE_Q_pipe_write_data(35 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_NUMBER_OF_SERVERS_1141_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NUMBER_OF_SERVERS_1141_inst_req_0;
      WPIPE_NUMBER_OF_SERVERS_1141_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NUMBER_OF_SERVERS_1141_inst_req_1;
      WPIPE_NUMBER_OF_SERVERS_1141_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_server_num_1118(0);
      data_in <= array_obj_ref_1143_wire;
      NUMBER_OF_SERVERS_write_3_gI: SplitGuardInterface generic map(name => "NUMBER_OF_SERVERS_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NUMBER_OF_SERVERS_write_3: OutputPortRevised -- 
        generic map ( name => "NUMBER_OF_SERVERS", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NUMBER_OF_SERVERS_pipe_write_req(0),
          oack => NUMBER_OF_SERVERS_pipe_write_ack(0),
          odata => NUMBER_OF_SERVERS_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared call operator group (0) : call_stmt_1219_call 
    UpdateRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(73 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1219_call_req_0;
      call_stmt_1219_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1219_call_req_1;
      call_stmt_1219_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not rwbar_1177_delayed_5_0_1203(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      UpdateRegister_call_group_0_gI: SplitGuardInterface generic map(name => "UpdateRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= bmask_1178_delayed_5_0_1206 & rval_1200 & wdata_1180_delayed_5_0_1209 & index_1181_delayed_5_0_1212;
      wval_1219 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 74,
        owidth => 74,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => UpdateRegister_call_reqs(0),
          ackR => UpdateRegister_call_acks(0),
          dataR => UpdateRegister_call_data(73 downto 0),
          tagR => UpdateRegister_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => UpdateRegister_return_acks(0), -- cross-over
          ackL => UpdateRegister_return_reqs(0), -- cross-over
          dataL => UpdateRegister_return_data(31 downto 0),
          tagL => UpdateRegister_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end SoftwareRegisterAccessDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity UpdateRegister is -- 
  generic (tag_length : integer); 
  port ( -- 
    bmask : in  std_logic_vector(3 downto 0);
    rval : in  std_logic_vector(31 downto 0);
    wdata : in  std_logic_vector(31 downto 0);
    index : in  std_logic_vector(5 downto 0);
    wval : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity UpdateRegister;
architecture UpdateRegister_arch of UpdateRegister is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 74)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal bmask_buffer :  std_logic_vector(3 downto 0);
  signal bmask_update_enable: Boolean;
  signal rval_buffer :  std_logic_vector(31 downto 0);
  signal rval_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(31 downto 0);
  signal wdata_update_enable: Boolean;
  signal index_buffer :  std_logic_vector(5 downto 0);
  signal index_update_enable: Boolean;
  -- output port buffer signals
  signal wval_buffer :  std_logic_vector(31 downto 0);
  signal wval_update_enable: Boolean;
  signal UpdateRegister_CP_34_start: Boolean;
  signal UpdateRegister_CP_34_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal CONCAT_u16_u32_170_inst_req_0 : boolean;
  signal CONCAT_u16_u32_170_inst_ack_0 : boolean;
  signal CONCAT_u16_u32_170_inst_req_1 : boolean;
  signal CONCAT_u16_u32_170_inst_ack_1 : boolean;
  signal array_obj_ref_173_store_0_req_0 : boolean;
  signal array_obj_ref_173_store_0_ack_0 : boolean;
  signal array_obj_ref_173_store_0_req_1 : boolean;
  signal array_obj_ref_173_store_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "UpdateRegister_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 74) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(3 downto 0) <= bmask;
  bmask_buffer <= in_buffer_data_out(3 downto 0);
  in_buffer_data_in(35 downto 4) <= rval;
  rval_buffer <= in_buffer_data_out(35 downto 4);
  in_buffer_data_in(67 downto 36) <= wdata;
  wdata_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(73 downto 68) <= index;
  index_buffer <= in_buffer_data_out(73 downto 68);
  in_buffer_data_in(tag_length + 73 downto 74) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 73 downto 74);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  UpdateRegister_CP_34_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "UpdateRegister_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= wval_buffer;
  wval <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= UpdateRegister_CP_34_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= UpdateRegister_CP_34_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= UpdateRegister_CP_34_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  UpdateRegister_CP_34: Block -- control-path 
    signal UpdateRegister_CP_34_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    UpdateRegister_CP_34_elements(0) <= UpdateRegister_CP_34_start;
    UpdateRegister_CP_34_symbol <= UpdateRegister_CP_34_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (39) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_sample_start_
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_update_start_
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Sample/rr
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Update/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Update/cr
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_update_start_
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_offset_calculated
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_resized_0
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_scaled_0
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_computed_0
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_resize_0/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_resize_0/$exit
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_resize_0/index_resize_req
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_resize_0/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_scale_0/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_scale_0/$exit
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_scale_0/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_scale_0/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_final_index_sum_regn/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_final_index_sum_regn/$exit
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_final_index_sum_regn/req
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_final_index_sum_regn/ack
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_base_plus_offset/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_base_plus_offset/$exit
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_word_addrgen/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_word_addrgen/$exit
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_word_addrgen/root_register_req
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_word_addrgen/root_register_ack
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/word_access_complete/word_0/cr
      -- 
    rr_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(0), ack => CONCAT_u16_u32_170_inst_req_0); -- 
    cr_52_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_52_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(0), ack => CONCAT_u16_u32_170_inst_req_1); -- 
    cr_114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(0), ack => array_obj_ref_173_store_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_sample_completed_
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Sample/ra
      -- 
    ra_48_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_170_inst_ack_0, ack => UpdateRegister_CP_34_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_update_completed_
      -- CP-element group 2: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Update/$exit
      -- CP-element group 2: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Update/ca
      -- 
    ca_53_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_170_inst_ack_1, ack => UpdateRegister_CP_34_elements(2)); -- 
    -- CP-element group 3:  join  transition  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_sample_start_
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/$entry
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/array_obj_ref_173_Split/$entry
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/array_obj_ref_173_Split/$exit
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/array_obj_ref_173_Split/split_req
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/array_obj_ref_173_Split/split_ack
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/word_access_start/$entry
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/word_access_start/word_0/rr
      -- 
    rr_103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(3), ack => array_obj_ref_173_store_0_req_0); -- 
    UpdateRegister_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "UpdateRegister_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= UpdateRegister_CP_34_elements(0) & UpdateRegister_CP_34_elements(2);
      gj_UpdateRegister_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => UpdateRegister_CP_34_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_sample_completed_
      -- CP-element group 4: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/$exit
      -- CP-element group 4: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/word_access_start/$exit
      -- CP-element group 4: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/word_access_start/word_0/$exit
      -- CP-element group 4: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/word_access_start/word_0/ra
      -- 
    ra_104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_173_store_0_ack_0, ack => UpdateRegister_CP_34_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (7) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_175/$exit
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_update_completed_
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/$exit
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/word_access_complete/$exit
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/word_access_complete/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/word_access_complete/word_0/ca
      -- 
    ca_115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_173_store_0_ack_1, ack => UpdateRegister_CP_34_elements(5)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u8_u16_160_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_169_wire : std_logic_vector(15 downto 0);
    signal MUX_155_wire : std_logic_vector(7 downto 0);
    signal MUX_159_wire : std_logic_vector(7 downto 0);
    signal MUX_164_wire : std_logic_vector(7 downto 0);
    signal MUX_168_wire : std_logic_vector(7 downto 0);
    signal R_index_172_resized : std_logic_vector(5 downto 0);
    signal R_index_172_scaled : std_logic_vector(5 downto 0);
    signal array_obj_ref_173_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_173_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_173_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_173_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_173_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_173_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_173_word_offset_0 : std_logic_vector(5 downto 0);
    signal b0_106 : std_logic_vector(0 downto 0);
    signal b1_110 : std_logic_vector(0 downto 0);
    signal b2_114 : std_logic_vector(0 downto 0);
    signal b3_118 : std_logic_vector(0 downto 0);
    signal r0_122 : std_logic_vector(7 downto 0);
    signal r1_126 : std_logic_vector(7 downto 0);
    signal r2_130 : std_logic_vector(7 downto 0);
    signal r3_134 : std_logic_vector(7 downto 0);
    signal w0_138 : std_logic_vector(7 downto 0);
    signal w1_142 : std_logic_vector(7 downto 0);
    signal w2_146 : std_logic_vector(7 downto 0);
    signal w3_150 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_173_offset_scale_factor_0 <= "000001";
    array_obj_ref_173_resized_base_address <= "000000";
    array_obj_ref_173_word_offset_0 <= "000000";
    -- flow-through select operator MUX_155_inst
    MUX_155_wire <= w0_138 when (b0_106(0) /=  '0') else r0_122;
    -- flow-through select operator MUX_159_inst
    MUX_159_wire <= w1_142 when (b1_110(0) /=  '0') else r1_126;
    -- flow-through select operator MUX_164_inst
    MUX_164_wire <= w2_146 when (b2_114(0) /=  '0') else r2_130;
    -- flow-through select operator MUX_168_inst
    MUX_168_wire <= w3_150 when (b3_118(0) /=  '0') else r3_134;
    -- flow-through slice operator slice_105_inst
    b0_106 <= bmask_buffer(3 downto 3);
    -- flow-through slice operator slice_109_inst
    b1_110 <= bmask_buffer(2 downto 2);
    -- flow-through slice operator slice_113_inst
    b2_114 <= bmask_buffer(1 downto 1);
    -- flow-through slice operator slice_117_inst
    b3_118 <= bmask_buffer(0 downto 0);
    -- flow-through slice operator slice_121_inst
    r0_122 <= rval_buffer(31 downto 24);
    -- flow-through slice operator slice_125_inst
    r1_126 <= rval_buffer(23 downto 16);
    -- flow-through slice operator slice_129_inst
    r2_130 <= rval_buffer(15 downto 8);
    -- flow-through slice operator slice_133_inst
    r3_134 <= rval_buffer(7 downto 0);
    -- flow-through slice operator slice_137_inst
    w0_138 <= wdata_buffer(31 downto 24);
    -- flow-through slice operator slice_141_inst
    w1_142 <= wdata_buffer(23 downto 16);
    -- flow-through slice operator slice_145_inst
    w2_146 <= wdata_buffer(15 downto 8);
    -- flow-through slice operator slice_149_inst
    w3_150 <= wdata_buffer(7 downto 0);
    -- equivalence array_obj_ref_173_addr_0
    process(array_obj_ref_173_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_173_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_173_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_173_gather_scatter
    process(wval_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := wval_buffer;
      ov(31 downto 0) := iv;
      array_obj_ref_173_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_173_index_0_rename
    process(R_index_172_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_172_resized;
      ov(5 downto 0) := iv;
      R_index_172_scaled <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_173_index_0_resize
    process(index_buffer) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_buffer;
      ov(5 downto 0) := iv;
      R_index_172_resized <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_173_index_offset
    process(R_index_172_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_172_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_173_final_offset <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_173_root_address_inst
    process(array_obj_ref_173_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_173_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_173_root_address <= ov(5 downto 0);
      --
    end process;
    -- shared split operator group (0) : CONCAT_u16_u32_170_inst 
    ApConcat_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u8_u16_160_wire & CONCAT_u8_u16_169_wire;
      wval_buffer <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u16_u32_170_inst_req_0;
      CONCAT_u16_u32_170_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u16_u32_170_inst_req_1;
      CONCAT_u16_u32_170_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_0_gI: SplitGuardInterface generic map(name => "ApConcat_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator CONCAT_u8_u16_160_inst
    process(MUX_155_wire, MUX_159_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_155_wire, MUX_159_wire, tmp_var);
      CONCAT_u8_u16_160_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_169_inst
    process(MUX_164_wire, MUX_168_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_164_wire, MUX_168_wire, tmp_var);
      CONCAT_u8_u16_169_wire <= tmp_var; --
    end process;
    -- shared store operator group (0) : array_obj_ref_173_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_173_store_0_req_0;
      array_obj_ref_173_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_173_store_0_req_1;
      array_obj_ref_173_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_173_word_address_0;
      data_in <= array_obj_ref_173_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 6,
        data_width => 32,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(5 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end UpdateRegister_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity accessMemory is -- 
  generic (tag_length : integer); 
  port ( -- 
    lock : in  std_logic_vector(0 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    bmask : in  std_logic_vector(7 downto 0);
    addr : in  std_logic_vector(35 downto 0);
    wdata : in  std_logic_vector(63 downto 0);
    rdata : out  std_logic_vector(63 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMemory;
architecture accessMemory_arch of accessMemory is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 110)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal bmask_buffer :  std_logic_vector(7 downto 0);
  signal bmask_update_enable: Boolean;
  signal addr_buffer :  std_logic_vector(35 downto 0);
  signal addr_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(63 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(63 downto 0);
  signal rdata_update_enable: Boolean;
  signal accessMemory_CP_329_start: Boolean;
  signal accessMemory_CP_329_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_req_0 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_ack_0 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_req_1 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_ack_1 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_req_0 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_ack_0 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_req_1 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMemory_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 110) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= lock;
  lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(1 downto 1) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(1 downto 1);
  in_buffer_data_in(9 downto 2) <= bmask;
  bmask_buffer <= in_buffer_data_out(9 downto 2);
  in_buffer_data_in(45 downto 10) <= addr;
  addr_buffer <= in_buffer_data_out(45 downto 10);
  in_buffer_data_in(109 downto 46) <= wdata;
  wdata_buffer <= in_buffer_data_out(109 downto 46);
  in_buffer_data_in(tag_length + 109 downto 110) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 109 downto 110);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1,6 => 15);
    constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1,6 => 15);
    constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 7); -- 
  begin -- 
    preds <= lock_update_enable & rwbar_update_enable & bmask_update_enable & addr_update_enable & wdata_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMemory_CP_329_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMemory_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemory_CP_329_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  rdata_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 24) := "rdata_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_rdata_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => rdata_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 15,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMemory_CP_329_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemory_CP_329_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMemory_CP_329: Block -- control-path 
    signal accessMemory_CP_329_elements: BooleanArray(22 downto 0);
    -- 
  begin -- 
    accessMemory_CP_329_elements(0) <= accessMemory_CP_329_start;
    accessMemory_CP_329_symbol <= accessMemory_CP_329_elements(22);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	8 
    -- CP-element group 1: 	11 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_267_to_stmt_287/$entry
      -- 
    accessMemory_CP_329_elements(1) <= accessMemory_CP_329_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	9 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	16 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_267_to_stmt_287/lock_update_enable
      -- CP-element group 2: 	 assign_stmt_267_to_stmt_287/lock_update_enable_out
      -- 
    accessMemory_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_329_elements(9);
      gj_accessMemory_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	9 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	17 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_267_to_stmt_287/rwbar_update_enable
      -- CP-element group 3: 	 assign_stmt_267_to_stmt_287/rwbar_update_enable_out
      -- 
    accessMemory_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_329_elements(9);
      gj_accessMemory_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	9 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	18 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_267_to_stmt_287/bmask_update_enable
      -- CP-element group 4: 	 assign_stmt_267_to_stmt_287/bmask_update_enable_out
      -- 
    accessMemory_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_329_elements(9);
      gj_accessMemory_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	9 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	19 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_267_to_stmt_287/addr_update_enable
      -- CP-element group 5: 	 assign_stmt_267_to_stmt_287/addr_update_enable_out
      -- 
    accessMemory_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_329_elements(9);
      gj_accessMemory_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	9 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	20 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 assign_stmt_267_to_stmt_287/wdata_update_enable
      -- CP-element group 6: 	 assign_stmt_267_to_stmt_287/wdata_update_enable_out
      -- 
    accessMemory_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_329_elements(9);
      gj_accessMemory_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	21 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	12 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_267_to_stmt_287/rdata_update_enable
      -- CP-element group 7: 	 assign_stmt_267_to_stmt_287/rdata_update_enable_in
      -- 
    accessMemory_CP_329_elements(7) <= accessMemory_CP_329_elements(21);
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	10 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_sample_start_
      -- CP-element group 8: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Sample/$entry
      -- CP-element group 8: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Sample/req
      -- 
    req_354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_329_elements(8), ack => WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_req_0); -- 
    accessMemory_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_329_elements(1) & accessMemory_CP_329_elements(10);
      gj_accessMemory_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: 	3 
    -- CP-element group 9: 	4 
    -- CP-element group 9: 	5 
    -- CP-element group 9: 	6 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_sample_completed_
      -- CP-element group 9: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_update_start_
      -- CP-element group 9: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Sample/$exit
      -- CP-element group 9: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Sample/ack
      -- CP-element group 9: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Update/$entry
      -- CP-element group 9: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Update/req
      -- 
    ack_355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_ack_0, ack => accessMemory_CP_329_elements(9)); -- 
    req_359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_329_elements(9), ack => WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: marked-successors 
    -- CP-element group 10: 	8 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_update_completed_
      -- CP-element group 10: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Update/$exit
      -- CP-element group 10: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Update/ack
      -- 
    ack_360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_ack_1, ack => accessMemory_CP_329_elements(10)); -- 
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	1 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_sample_start_
      -- CP-element group 11: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Sample/$entry
      -- CP-element group 11: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Sample/rr
      -- 
    rr_368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_329_elements(11), ack => RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_req_0); -- 
    accessMemory_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessMemory_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_329_elements(1) & accessMemory_CP_329_elements(14);
      gj_accessMemory_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	7 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_update_start_
      -- CP-element group 12: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Update/$entry
      -- CP-element group 12: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Update/cr
      -- 
    cr_373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_329_elements(12), ack => RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_req_1); -- 
    accessMemory_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessMemory_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_329_elements(13) & accessMemory_CP_329_elements(7);
      gj_accessMemory_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	12 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_sample_completed_
      -- CP-element group 13: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Sample/$exit
      -- CP-element group 13: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Sample/ra
      -- 
    ra_369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_ack_0, ack => accessMemory_CP_329_elements(13)); -- 
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_update_completed_
      -- CP-element group 14: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Update/$exit
      -- CP-element group 14: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Update/ca
      -- 
    ca_374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_ack_1, ack => accessMemory_CP_329_elements(14)); -- 
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	22 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 assign_stmt_267_to_stmt_287/$exit
      -- 
    accessMemory_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessMemory_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_329_elements(14) & accessMemory_CP_329_elements(10);
      gj_accessMemory_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 lock_update_enable
      -- 
    accessMemory_CP_329_elements(16) <= accessMemory_CP_329_elements(2);
    -- CP-element group 17:  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	3 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 rwbar_update_enable
      -- 
    accessMemory_CP_329_elements(17) <= accessMemory_CP_329_elements(3);
    -- CP-element group 18:  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	4 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 bmask_update_enable
      -- 
    accessMemory_CP_329_elements(18) <= accessMemory_CP_329_elements(4);
    -- CP-element group 19:  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	5 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 addr_update_enable
      -- 
    accessMemory_CP_329_elements(19) <= accessMemory_CP_329_elements(5);
    -- CP-element group 20:  place  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	6 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 wdata_update_enable
      -- 
    accessMemory_CP_329_elements(20) <= accessMemory_CP_329_elements(6);
    -- CP-element group 21:  place  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	7 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 rdata_update_enable
      -- 
    -- CP-element group 22:  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 $exit
      -- 
    accessMemory_CP_329_elements(22) <= accessMemory_CP_329_elements(15);
    --  hookup: inputs to control-path 
    accessMemory_CP_329_elements(21) <= rdata_update_enable;
    -- hookup: output from control-path 
    lock_update_enable <= accessMemory_CP_329_elements(16);
    rwbar_update_enable <= accessMemory_CP_329_elements(17);
    bmask_update_enable <= accessMemory_CP_329_elements(18);
    addr_update_enable <= accessMemory_CP_329_elements(19);
    wdata_update_enable <= accessMemory_CP_329_elements(20);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u2_260_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u10_262_wire : std_logic_vector(9 downto 0);
    signal CONCAT_u36_u100_265_wire : std_logic_vector(99 downto 0);
    signal err_277 : std_logic_vector(0 downto 0);
    signal request_267 : std_logic_vector(109 downto 0);
    signal response_273 : std_logic_vector(64 downto 0);
    -- 
  begin -- 
    -- flow-through slice operator slice_276_inst
    err_277 <= response_273(64 downto 64);
    -- flow-through slice operator slice_280_inst
    rdata_buffer <= response_273(63 downto 0);
    -- binary operator CONCAT_u10_u110_266_inst
    process(CONCAT_u2_u10_262_wire, CONCAT_u36_u100_265_wire) -- 
      variable tmp_var : std_logic_vector(109 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u10_262_wire, CONCAT_u36_u100_265_wire, tmp_var);
      request_267 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_260_inst
    process(lock_buffer, rwbar_buffer) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(lock_buffer, rwbar_buffer, tmp_var);
      CONCAT_u1_u2_260_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u10_262_inst
    process(CONCAT_u1_u2_260_wire, bmask_buffer) -- 
      variable tmp_var : std_logic_vector(9 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_260_wire, bmask_buffer, tmp_var);
      CONCAT_u2_u10_262_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u36_u100_265_inst
    process(addr_buffer, wdata_buffer) -- 
      variable tmp_var : std_logic_vector(99 downto 0); -- 
    begin -- 
      ApConcat_proc(addr_buffer, wdata_buffer, tmp_var);
      CONCAT_u36_u100_265_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(64 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_req_0;
      RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_req_1;
      RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      response_273 <= data_out(64 downto 0);
      MEMORY_TO_NIC_RESPONSE_read_0_gI: SplitGuardInterface generic map(name => "MEMORY_TO_NIC_RESPONSE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      MEMORY_TO_NIC_RESPONSE_read_0: InputPortRevised -- 
        generic map ( name => "MEMORY_TO_NIC_RESPONSE_read_0", data_width => 65,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => MEMORY_TO_NIC_RESPONSE_pipe_read_req(0),
          oack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack(0),
          odata => MEMORY_TO_NIC_RESPONSE_pipe_read_data(64 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_NIC_TO_MEMORY_REQUEST_268_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_req_0;
      WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_req_1;
      WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= request_267;
      NIC_TO_MEMORY_REQUEST_write_0_gI: SplitGuardInterface generic map(name => "NIC_TO_MEMORY_REQUEST_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_TO_MEMORY_REQUEST_write_0: OutputPortRevised -- 
        generic map ( name => "NIC_TO_MEMORY_REQUEST", data_width => 110, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_TO_MEMORY_REQUEST_pipe_write_req(0),
          oack => NIC_TO_MEMORY_REQUEST_pipe_write_ack(0),
          odata => NIC_TO_MEMORY_REQUEST_pipe_write_data(109 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end accessMemory_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity acquireMutex is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    m_ok : out  std_logic_vector(0 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity acquireMutex;
architecture acquireMutex_arch of acquireMutex is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal m_ok_buffer :  std_logic_vector(0 downto 0);
  signal acquireMutex_CP_381_start: Boolean;
  signal acquireMutex_CP_381_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal if_stmt_313_branch_ack_0 : boolean;
  signal call_stmt_308_call_req_1 : boolean;
  signal if_stmt_313_branch_ack_1 : boolean;
  signal if_stmt_313_branch_req_0 : boolean;
  signal call_stmt_327_call_ack_1 : boolean;
  signal call_stmt_327_call_req_1 : boolean;
  signal call_stmt_327_call_ack_0 : boolean;
  signal call_stmt_327_call_req_0 : boolean;
  signal call_stmt_308_call_ack_0 : boolean;
  signal call_stmt_347_call_ack_1 : boolean;
  signal call_stmt_347_call_req_1 : boolean;
  signal call_stmt_308_call_req_0 : boolean;
  signal call_stmt_347_call_ack_0 : boolean;
  signal call_stmt_347_call_req_0 : boolean;
  signal call_stmt_308_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "acquireMutex_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  acquireMutex_CP_381_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "acquireMutex_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  m_ok_buffer <= "1";
  out_buffer_data_in(0 downto 0) <= m_ok_buffer;
  m_ok <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= acquireMutex_CP_381_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= acquireMutex_CP_381_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= acquireMutex_CP_381_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  acquireMutex_CP_381: Block -- control-path 
    signal acquireMutex_CP_381_elements: BooleanArray(9 downto 0);
    -- 
  begin -- 
    acquireMutex_CP_381_elements(0) <= acquireMutex_CP_381_start;
    acquireMutex_CP_381_symbol <= acquireMutex_CP_381_elements(8);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	9 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 branch_block_stmt_292/assign_stmt_295/$exit
      -- CP-element group 0: 	 branch_block_stmt_292/assign_stmt_295/$entry
      -- CP-element group 0: 	 branch_block_stmt_292/merge_stmt_296__entry___PhiReq/$exit
      -- CP-element group 0: 	 branch_block_stmt_292/merge_stmt_296__entry__
      -- CP-element group 0: 	 branch_block_stmt_292/merge_stmt_296__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_292/assign_stmt_295__exit__
      -- CP-element group 0: 	 branch_block_stmt_292/assign_stmt_295__entry__
      -- CP-element group 0: 	 branch_block_stmt_292/merge_stmt_296_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_292/branch_block_stmt_292__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_292/$entry
      -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	9 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_Sample/cra
      -- CP-element group 1: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_sample_completed_
      -- 
    cra_413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_308_call_ack_0, ack => acquireMutex_CP_381_elements(1)); -- 
    -- CP-element group 2:  branch  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	9 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (27) 
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_else_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312__exit__
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_if_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/EQ_u32_u1_316_place
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/branch_req
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/$exit
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/EQ_u32_u1_316_inputs/$exit
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/$exit
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/Update/ca
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/EQ_u32_u1_316_inputs/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/$exit
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/Update/cr
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/$exit
      -- CP-element group 2: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313__entry__
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_Update/cca
      -- 
    cca_418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_308_call_ack_1, ack => acquireMutex_CP_381_elements(2)); -- 
    branch_req_445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireMutex_CP_381_elements(2), ack => if_stmt_313_branch_req_0); -- 
    -- CP-element group 3:  fork  transition  place  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	5 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (10) 
      -- CP-element group 3: 	 branch_block_stmt_292/if_stmt_313_if_link/if_choice_transition
      -- CP-element group 3: 	 branch_block_stmt_292/if_stmt_313_if_link/$exit
      -- CP-element group 3: 	 branch_block_stmt_292/call_stmt_327/call_stmt_327_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_292/call_stmt_327/call_stmt_327_Update/ccr
      -- CP-element group 3: 	 branch_block_stmt_292/call_stmt_327/call_stmt_327_Sample/crr
      -- CP-element group 3: 	 branch_block_stmt_292/call_stmt_327/call_stmt_327_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_292/call_stmt_327/call_stmt_327_update_start_
      -- CP-element group 3: 	 branch_block_stmt_292/call_stmt_327/call_stmt_327_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_292/call_stmt_327/$entry
      -- CP-element group 3: 	 branch_block_stmt_292/call_stmt_327__entry__
      -- 
    if_choice_transition_450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_313_branch_ack_1, ack => acquireMutex_CP_381_elements(3)); -- 
    ccr_473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireMutex_CP_381_elements(3), ack => call_stmt_327_call_req_1); -- 
    crr_468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireMutex_CP_381_elements(3), ack => call_stmt_327_call_req_0); -- 
    -- CP-element group 4:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4: 	8 
    -- CP-element group 4:  members (11) 
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_313_else_link/$exit
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_313_else_link/else_choice_transition
      -- CP-element group 4: 	 branch_block_stmt_292/assign_stmt_336_to_call_stmt_347/$entry
      -- CP-element group 4: 	 branch_block_stmt_292/assign_stmt_336_to_call_stmt_347/call_stmt_347_Update/ccr
      -- CP-element group 4: 	 branch_block_stmt_292/assign_stmt_336_to_call_stmt_347/call_stmt_347_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_292/assign_stmt_336_to_call_stmt_347/call_stmt_347_Sample/crr
      -- CP-element group 4: 	 branch_block_stmt_292/assign_stmt_336_to_call_stmt_347/call_stmt_347_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_292/assign_stmt_336_to_call_stmt_347/call_stmt_347_update_start_
      -- CP-element group 4: 	 branch_block_stmt_292/assign_stmt_336_to_call_stmt_347__entry__
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_313__exit__
      -- CP-element group 4: 	 branch_block_stmt_292/assign_stmt_336_to_call_stmt_347/call_stmt_347_sample_start_
      -- 
    else_choice_transition_454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_313_branch_ack_0, ack => acquireMutex_CP_381_elements(4)); -- 
    ccr_490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireMutex_CP_381_elements(4), ack => call_stmt_347_call_req_1); -- 
    crr_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireMutex_CP_381_elements(4), ack => call_stmt_347_call_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	3 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_292/call_stmt_327/call_stmt_327_Sample/cra
      -- CP-element group 5: 	 branch_block_stmt_292/call_stmt_327/call_stmt_327_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_292/call_stmt_327/call_stmt_327_sample_completed_
      -- 
    cra_469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_327_call_ack_0, ack => acquireMutex_CP_381_elements(5)); -- 
    -- CP-element group 6:  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (8) 
      -- CP-element group 6: 	 branch_block_stmt_292/call_stmt_327/call_stmt_327_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_292/call_stmt_327/call_stmt_327_Update/cca
      -- CP-element group 6: 	 branch_block_stmt_292/loopback_PhiReq/$exit
      -- CP-element group 6: 	 branch_block_stmt_292/loopback_PhiReq/$entry
      -- CP-element group 6: 	 branch_block_stmt_292/call_stmt_327/call_stmt_327_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_292/call_stmt_327/$exit
      -- CP-element group 6: 	 branch_block_stmt_292/loopback
      -- CP-element group 6: 	 branch_block_stmt_292/call_stmt_327__exit__
      -- 
    cca_474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_327_call_ack_1, ack => acquireMutex_CP_381_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_292/assign_stmt_336_to_call_stmt_347/call_stmt_347_Sample/cra
      -- CP-element group 7: 	 branch_block_stmt_292/assign_stmt_336_to_call_stmt_347/call_stmt_347_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_292/assign_stmt_336_to_call_stmt_347/call_stmt_347_sample_completed_
      -- 
    cra_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_347_call_ack_0, ack => acquireMutex_CP_381_elements(7)); -- 
    -- CP-element group 8:  transition  place  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	4 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (10) 
      -- CP-element group 8: 	 $exit
      -- CP-element group 8: 	 branch_block_stmt_292/assign_stmt_336_to_call_stmt_347/call_stmt_347_Update/cca
      -- CP-element group 8: 	 branch_block_stmt_292/assign_stmt_336_to_call_stmt_347/call_stmt_347_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_292/branch_block_stmt_292__exit__
      -- CP-element group 8: 	 branch_block_stmt_292/assign_stmt_336_to_call_stmt_347/call_stmt_347_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_292/assign_stmt_336_to_call_stmt_347__exit__
      -- CP-element group 8: 	 branch_block_stmt_292/$exit
      -- CP-element group 8: 	 assign_stmt_352/$exit
      -- CP-element group 8: 	 assign_stmt_352/$entry
      -- CP-element group 8: 	 branch_block_stmt_292/assign_stmt_336_to_call_stmt_347/$exit
      -- 
    cca_491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_347_call_ack_1, ack => acquireMutex_CP_381_elements(8)); -- 
    -- CP-element group 9:  merge  fork  transition  place  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: 	2 
    -- CP-element group 9:  members (13) 
      -- CP-element group 9: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_Update/ccr
      -- CP-element group 9: 	 branch_block_stmt_292/merge_stmt_296_PhiAck/dummy
      -- CP-element group 9: 	 branch_block_stmt_292/merge_stmt_296_PhiAck/$exit
      -- CP-element group 9: 	 branch_block_stmt_292/merge_stmt_296_PhiAck/$entry
      -- CP-element group 9: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312__entry__
      -- CP-element group 9: 	 branch_block_stmt_292/merge_stmt_296_PhiReqMerge
      -- CP-element group 9: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/$entry
      -- CP-element group 9: 	 branch_block_stmt_292/merge_stmt_296__exit__
      -- CP-element group 9: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_Sample/crr
      -- CP-element group 9: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_update_start_
      -- CP-element group 9: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_sample_start_
      -- 
    ccr_417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireMutex_CP_381_elements(9), ack => call_stmt_308_call_req_1); -- 
    crr_412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireMutex_CP_381_elements(9), ack => call_stmt_308_call_req_0); -- 
    acquireMutex_CP_381_elements(9) <= OrReduce(acquireMutex_CP_381_elements(0) & acquireMutex_CP_381_elements(6));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u32_u1_316_wire : std_logic_vector(0 downto 0);
    signal NOT_u8_u8_303_wire_constant : std_logic_vector(7 downto 0);
    signal NOT_u8_u8_323_wire_constant : std_logic_vector(7 downto 0);
    signal NOT_u8_u8_343_wire_constant : std_logic_vector(7 downto 0);
    signal err_327 : std_logic_vector(63 downto 0);
    signal ignore_347 : std_logic_vector(63 downto 0);
    signal konst_315_wire_constant : std_logic_vector(31 downto 0);
    signal mutex_address_295 : std_logic_vector(35 downto 0);
    signal mutex_plus_nentries_308 : std_logic_vector(63 downto 0);
    signal mutex_val_312 : std_logic_vector(31 downto 0);
    signal slice_334_wire : std_logic_vector(31 downto 0);
    signal type_cast_298_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_300_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_306_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_318_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_320_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_332_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_338_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_340_wire_constant : std_logic_vector(0 downto 0);
    signal wval_336 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_303_wire_constant <= "11111111";
    NOT_u8_u8_323_wire_constant <= "11111111";
    NOT_u8_u8_343_wire_constant <= "11111111";
    konst_315_wire_constant <= "00000000000000000000000000000001";
    type_cast_298_wire_constant <= "1";
    type_cast_300_wire_constant <= "1";
    type_cast_306_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_318_wire_constant <= "0";
    type_cast_320_wire_constant <= "1";
    type_cast_332_wire_constant <= "00000000000000000000000000000001";
    type_cast_338_wire_constant <= "0";
    type_cast_340_wire_constant <= "0";
    -- flow-through slice operator slice_311_inst
    mutex_val_312 <= mutex_plus_nentries_308(63 downto 32);
    -- flow-through slice operator slice_334_inst
    slice_334_wire <= mutex_plus_nentries_308(31 downto 0);
    -- interlock W_mutex_address_293_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 35 downto 0) := q_base_address_buffer(35 downto 0);
      mutex_address_295 <= tmp_var; -- 
    end process;
    if_stmt_313_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u32_u1_316_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_313_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_313_branch_req_0,
          ack0 => if_stmt_313_branch_ack_0,
          ack1 => if_stmt_313_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u32_u64_335_inst
    process(type_cast_332_wire_constant, slice_334_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_332_wire_constant, slice_334_wire, tmp_var);
      wval_336 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_316_inst
    process(mutex_val_312) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(mutex_val_312, konst_315_wire_constant, tmp_var);
      EQ_u32_u1_316_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_327_call call_stmt_308_call call_stmt_347_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(329 downto 0);
      signal data_out: std_logic_vector(191 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= call_stmt_327_call_req_0;
      reqL_unguarded(1) <= call_stmt_308_call_req_0;
      reqL_unguarded(0) <= call_stmt_347_call_req_0;
      call_stmt_327_call_ack_0 <= ackL_unguarded(2);
      call_stmt_308_call_ack_0 <= ackL_unguarded(1);
      call_stmt_347_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= call_stmt_327_call_req_1;
      reqR_unguarded(1) <= call_stmt_308_call_req_1;
      reqR_unguarded(0) <= call_stmt_347_call_req_1;
      call_stmt_327_call_ack_1 <= ackR_unguarded(2);
      call_stmt_308_call_ack_1 <= ackR_unguarded(1);
      call_stmt_347_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_2: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_318_wire_constant & type_cast_320_wire_constant & NOT_u8_u8_323_wire_constant & mutex_address_295 & mutex_plus_nentries_308 & type_cast_298_wire_constant & type_cast_300_wire_constant & NOT_u8_u8_303_wire_constant & mutex_address_295 & type_cast_306_wire_constant & type_cast_338_wire_constant & type_cast_340_wire_constant & NOT_u8_u8_343_wire_constant & mutex_address_295 & wval_336;
      err_327 <= data_out(191 downto 128);
      mutex_plus_nentries_308 <= data_out(127 downto 64);
      ignore_347 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 330,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 3,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 192,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 3) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end acquireMutex_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity delay_time_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    T : in  std_logic_vector(31 downto 0);
    delay_done : out  std_logic_vector(0 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity delay_time_Operator;
architecture delay_time_Operator_arch of delay_time_Operator is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal update_ack_symbol: Boolean;
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal T_buffer :  std_logic_vector(31 downto 0);
  signal T_update_enable: Boolean;
  signal T_update_enable_unmarked: Boolean;
  -- output port buffer signals
  signal delay_done_buffer :  std_logic_vector(0 downto 0);
  signal delay_time_CP_1231_start: Boolean;
  signal delay_time_CP_1231_symbol: Boolean;
  signal cp_all_inputs_sampled: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_856_branch_ack_1 : boolean;
  signal do_while_stmt_856_branch_ack_0 : boolean;
  signal do_while_stmt_856_branch_req_0 : boolean;
  signal phi_stmt_858_req_0 : boolean;
  signal phi_stmt_858_req_1 : boolean;
  signal phi_stmt_858_ack_0 : boolean;
  signal nR_867_860_buf_req_0 : boolean;
  signal nR_867_860_buf_ack_0 : boolean;
  signal nR_867_860_buf_req_1 : boolean;
  signal nR_867_860_buf_ack_1 : boolean;
  signal T_861_buf_req_0 : boolean;
  signal T_861_buf_ack_0 : boolean;
  signal T_861_buf_req_1 : boolean;
  signal T_861_buf_ack_1 : boolean;
  -- 
begin --  
  sample_ack <= delay_time_CP_1231_symbol;
  -- input handling ------------------------------------------------
  T_buffer <= T;
  delay_time_CP_1231_start <= sample_req;
  -- output handling  -------------------------------------------------------
  delay_done_buffer <= "1";
  delay_done <= delay_done_buffer;
  update_ack_symbol <= delay_time_CP_1231_symbol;
  update_ack <= update_ack_symbol;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  delay_time_CP_1231: Block -- control-path 
    signal delay_time_CP_1231_elements: BooleanArray(32 downto 0);
    -- 
  begin -- 
    delay_time_CP_1231_elements(0) <= delay_time_CP_1231_start;
    delay_time_CP_1231_symbol <= delay_time_CP_1231_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_855/$entry
      -- CP-element group 0: 	 branch_block_stmt_855/branch_block_stmt_855__entry__
      -- CP-element group 0: 	 branch_block_stmt_855/do_while_stmt_856__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	32 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (8) 
      -- CP-element group 1: 	 branch_block_stmt_855/assign_stmt_874/$exit
      -- CP-element group 1: 	 branch_block_stmt_855/assign_stmt_874/$entry
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_855/$exit
      -- CP-element group 1: 	 branch_block_stmt_855/branch_block_stmt_855__exit__
      -- CP-element group 1: 	 branch_block_stmt_855/do_while_stmt_856__exit__
      -- CP-element group 1: 	 branch_block_stmt_855/assign_stmt_874__entry__
      -- CP-element group 1: 	 branch_block_stmt_855/assign_stmt_874__exit__
      -- 
    delay_time_CP_1231_elements(1) <= delay_time_CP_1231_elements(32);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_855/do_while_stmt_856/$entry
      -- CP-element group 2: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856__entry__
      -- 
    delay_time_CP_1231_elements(2) <= delay_time_CP_1231_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	32 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856__exit__
      -- 
    -- Element group delay_time_CP_1231_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_855/do_while_stmt_856/loop_back
      -- 
    -- Element group delay_time_CP_1231_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	30 
    -- CP-element group 5: 	31 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_855/do_while_stmt_856/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_855/do_while_stmt_856/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_855/do_while_stmt_856/condition_done
      -- 
    delay_time_CP_1231_elements(5) <= delay_time_CP_1231_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	14 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_855/do_while_stmt_856/loop_body_done
      -- 
    delay_time_CP_1231_elements(6) <= delay_time_CP_1231_elements(14);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/back_edge_to_loop_body
      -- 
    delay_time_CP_1231_elements(7) <= delay_time_CP_1231_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/first_time_through_loop_body
      -- 
    delay_time_CP_1231_elements(8) <= delay_time_CP_1231_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	29 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/loop_body_start
      -- 
    -- Element group delay_time_CP_1231_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	29 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/condition_evaluated
      -- 
    condition_evaluated_1257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1231_elements(10), ack => do_while_stmt_856_branch_req_0); -- 
    delay_time_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1231_elements(15) & delay_time_CP_1231_elements(29);
      gj_delay_time_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1231_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/phi_stmt_858_sample_start__ps
      -- 
    delay_time_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1231_elements(12) & delay_time_CP_1231_elements(15);
      gj_delay_time_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1231_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/phi_stmt_858_sample_start_
      -- 
    delay_time_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1231_elements(9) & delay_time_CP_1231_elements(14);
      gj_delay_time_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1231_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/phi_stmt_858_update_start_
      -- CP-element group 13: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/phi_stmt_858_update_start__ps
      -- 
    delay_time_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1231_elements(9) & delay_time_CP_1231_elements(15);
      gj_delay_time_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1231_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	6 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (4) 
      -- CP-element group 14: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/$exit
      -- CP-element group 14: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/phi_stmt_858_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/phi_stmt_858_sample_completed__ps
      -- 
    -- Element group delay_time_CP_1231_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15: 	13 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/phi_stmt_858_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/phi_stmt_858_update_completed__ps
      -- 
    -- Element group delay_time_CP_1231_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/phi_stmt_858_loopback_trigger
      -- 
    delay_time_CP_1231_elements(16) <= delay_time_CP_1231_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/phi_stmt_858_loopback_sample_req
      -- CP-element group 17: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/phi_stmt_858_loopback_sample_req_ps
      -- 
    phi_stmt_858_loopback_sample_req_1272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_858_loopback_sample_req_1272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1231_elements(17), ack => phi_stmt_858_req_0); -- 
    -- Element group delay_time_CP_1231_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/phi_stmt_858_entry_trigger
      -- 
    delay_time_CP_1231_elements(18) <= delay_time_CP_1231_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/phi_stmt_858_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/phi_stmt_858_entry_sample_req_ps
      -- 
    phi_stmt_858_entry_sample_req_1275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_858_entry_sample_req_1275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1231_elements(19), ack => phi_stmt_858_req_1); -- 
    -- Element group delay_time_CP_1231_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/phi_stmt_858_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/phi_stmt_858_phi_mux_ack_ps
      -- 
    phi_stmt_858_phi_mux_ack_1278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_858_ack_0, ack => delay_time_CP_1231_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_nR_860_sample_start__ps
      -- CP-element group 21: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_nR_860_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_nR_860_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_nR_860_Sample/req
      -- 
    req_1291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1231_elements(21), ack => nR_867_860_buf_req_0); -- 
    -- Element group delay_time_CP_1231_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (4) 
      -- CP-element group 22: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_nR_860_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_nR_860_update_start_
      -- CP-element group 22: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_nR_860_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_nR_860_Update/req
      -- 
    req_1296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1231_elements(22), ack => nR_867_860_buf_req_1); -- 
    -- Element group delay_time_CP_1231_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (4) 
      -- CP-element group 23: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_nR_860_sample_completed__ps
      -- CP-element group 23: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_nR_860_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_nR_860_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_nR_860_Sample/ack
      -- 
    ack_1292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nR_867_860_buf_ack_0, ack => delay_time_CP_1231_elements(23)); -- 
    -- CP-element group 24:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_nR_860_update_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_nR_860_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_nR_860_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_nR_860_Update/ack
      -- 
    ack_1297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nR_867_860_buf_ack_1, ack => delay_time_CP_1231_elements(24)); -- 
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_T_861_sample_start__ps
      -- CP-element group 25: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_T_861_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_T_861_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_T_861_Sample/req
      -- 
    req_1309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1231_elements(25), ack => T_861_buf_req_0); -- 
    -- Element group delay_time_CP_1231_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_T_861_update_start__ps
      -- CP-element group 26: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_T_861_update_start_
      -- CP-element group 26: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_T_861_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_T_861_Update/req
      -- 
    req_1314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1231_elements(26), ack => T_861_buf_req_1); -- 
    -- Element group delay_time_CP_1231_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_T_861_sample_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_T_861_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_T_861_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_T_861_Sample/ack
      -- 
    ack_1310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => T_861_buf_ack_0, ack => delay_time_CP_1231_elements(27)); -- 
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_T_861_update_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_T_861_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_T_861_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/R_T_861_Update/ack
      -- 
    ack_1315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => T_861_buf_ack_1, ack => delay_time_CP_1231_elements(28)); -- 
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	9 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	10 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_855/do_while_stmt_856/do_while_stmt_856_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group delay_time_CP_1231_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => delay_time_CP_1231_elements(9), ack => delay_time_CP_1231_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	5 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_855/do_while_stmt_856/loop_exit/ack
      -- CP-element group 30: 	 branch_block_stmt_855/do_while_stmt_856/loop_exit/$exit
      -- 
    ack_1321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_856_branch_ack_0, ack => delay_time_CP_1231_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	5 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_855/do_while_stmt_856/loop_taken/ack
      -- CP-element group 31: 	 branch_block_stmt_855/do_while_stmt_856/loop_taken/$exit
      -- 
    ack_1325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_856_branch_ack_1, ack => delay_time_CP_1231_elements(31)); -- 
    -- CP-element group 32:  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	3 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	1 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_855/do_while_stmt_856/$exit
      -- 
    delay_time_CP_1231_elements(32) <= delay_time_CP_1231_elements(3);
    delay_time_do_while_stmt_856_terminator_1326: loop_terminator -- 
      generic map (name => " delay_time_do_while_stmt_856_terminator_1326", max_iterations_in_flight =>7) 
      port map(loop_body_exit => delay_time_CP_1231_elements(6),loop_continue => delay_time_CP_1231_elements(31),loop_terminate => delay_time_CP_1231_elements(30),loop_back => delay_time_CP_1231_elements(4),loop_exit => delay_time_CP_1231_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_858_phi_seq_1316_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= delay_time_CP_1231_elements(16);
      delay_time_CP_1231_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= delay_time_CP_1231_elements(23);
      delay_time_CP_1231_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= delay_time_CP_1231_elements(24);
      delay_time_CP_1231_elements(17) <= phi_mux_reqs(0);
      triggers(1)  <= delay_time_CP_1231_elements(18);
      delay_time_CP_1231_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= delay_time_CP_1231_elements(27);
      delay_time_CP_1231_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= delay_time_CP_1231_elements(28);
      delay_time_CP_1231_elements(19) <= phi_mux_reqs(1);
      phi_stmt_858_phi_seq_1316 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_858_phi_seq_1316") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => delay_time_CP_1231_elements(11), 
          phi_sample_ack => delay_time_CP_1231_elements(14), 
          phi_update_req => delay_time_CP_1231_elements(13), 
          phi_update_ack => delay_time_CP_1231_elements(15), 
          phi_mux_ack => delay_time_CP_1231_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1258_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= delay_time_CP_1231_elements(7);
        preds(1)  <= delay_time_CP_1231_elements(8);
        entry_tmerge_1258 : transition_merge -- 
          generic map(name => " entry_tmerge_1258")
          port map (preds => preds, symbol_out => delay_time_CP_1231_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_858 : std_logic_vector(31 downto 0);
    signal T_861_buffered : std_logic_vector(31 downto 0);
    signal UGT_u32_u1_871_wire : std_logic_vector(0 downto 0);
    signal konst_865_wire_constant : std_logic_vector(31 downto 0);
    signal konst_870_wire_constant : std_logic_vector(31 downto 0);
    signal nR_867 : std_logic_vector(31 downto 0);
    signal nR_867_860_buffered : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_865_wire_constant <= "00000000000000000000000000000001";
    konst_870_wire_constant <= "00000000000000000000000000000000";
    phi_stmt_858: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nR_867_860_buffered & T_861_buffered;
      req <= phi_stmt_858_req_0 & phi_stmt_858_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_858",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_858_ack_0,
          idata => idata,
          odata => R_858,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_858
    T_861_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= T_861_buf_req_0;
      T_861_buf_ack_0<= wack(0);
      rreq(0) <= T_861_buf_req_1;
      T_861_buf_ack_1<= rack(0);
      T_861_buf : InterlockBuffer generic map ( -- 
        name => "T_861_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => T_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => T_861_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nR_867_860_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nR_867_860_buf_req_0;
      nR_867_860_buf_ack_0<= wack(0);
      rreq(0) <= nR_867_860_buf_req_1;
      nR_867_860_buf_ack_1<= rack(0);
      nR_867_860_buf : InterlockBuffer generic map ( -- 
        name => "nR_867_860_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nR_867,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nR_867_860_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_856_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= UGT_u32_u1_871_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_856_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_856_branch_req_0,
          ack0 => do_while_stmt_856_branch_ack_0,
          ack1 => do_while_stmt_856_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator SUB_u32_u32_866_inst
    process(R_858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(R_858, konst_865_wire_constant, tmp_var);
      nR_867 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_871_inst
    process(R_858) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(R_858, konst_870_wire_constant, tmp_var);
      UGT_u32_u1_871_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end delay_time_Operator_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity getQueueElement is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    read_pointer : in  std_logic_vector(31 downto 0);
    q_r_data : out  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueueElement;
architecture getQueueElement_arch of getQueueElement is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 68)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal read_pointer_buffer :  std_logic_vector(31 downto 0);
  signal read_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal q_r_data_buffer :  std_logic_vector(31 downto 0);
  signal q_r_data_update_enable: Boolean;
  signal getQueueElement_CP_530_start: Boolean;
  signal getQueueElement_CP_530_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal MUX_434_inst_ack_0 : boolean;
  signal call_stmt_419_call_ack_0 : boolean;
  signal MUX_434_inst_req_0 : boolean;
  signal call_stmt_419_call_req_0 : boolean;
  signal MUX_434_inst_ack_1 : boolean;
  signal MUX_434_inst_req_1 : boolean;
  signal call_stmt_419_call_ack_1 : boolean;
  signal call_stmt_419_call_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueueElement_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 68) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= read_pointer;
  read_pointer_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(tag_length + 67 downto 68) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 67 downto 68);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueueElement_CP_530_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueueElement_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= q_r_data_buffer;
  q_r_data <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueElement_CP_530_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueueElement_CP_530_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueElement_CP_530_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueueElement_CP_530: Block -- control-path 
    signal getQueueElement_CP_530_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    getQueueElement_CP_530_elements(0) <= getQueueElement_CP_530_start;
    getQueueElement_CP_530_symbol <= getQueueElement_CP_530_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 assign_stmt_394_to_assign_stmt_435/call_stmt_419_Sample/crr
      -- CP-element group 0: 	 assign_stmt_394_to_assign_stmt_435/MUX_434_complete/$entry
      -- CP-element group 0: 	 assign_stmt_394_to_assign_stmt_435/MUX_434_complete/req
      -- CP-element group 0: 	 assign_stmt_394_to_assign_stmt_435/MUX_434_update_start_
      -- CP-element group 0: 	 assign_stmt_394_to_assign_stmt_435/call_stmt_419_sample_start_
      -- CP-element group 0: 	 assign_stmt_394_to_assign_stmt_435/call_stmt_419_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_394_to_assign_stmt_435/call_stmt_419_update_start_
      -- CP-element group 0: 	 assign_stmt_394_to_assign_stmt_435/call_stmt_419_Update/ccr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_394_to_assign_stmt_435/call_stmt_419_Update/$entry
      -- CP-element group 0: 	 assign_stmt_394_to_assign_stmt_435/$entry
      -- 
    crr_543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_530_elements(0), ack => call_stmt_419_call_req_0); -- 
    req_562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_530_elements(0), ack => MUX_434_inst_req_1); -- 
    ccr_548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_530_elements(0), ack => call_stmt_419_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_394_to_assign_stmt_435/call_stmt_419_Sample/cra
      -- CP-element group 1: 	 assign_stmt_394_to_assign_stmt_435/call_stmt_419_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_394_to_assign_stmt_435/call_stmt_419_sample_completed_
      -- 
    cra_544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_419_call_ack_0, ack => getQueueElement_CP_530_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_394_to_assign_stmt_435/MUX_434_start/$entry
      -- CP-element group 2: 	 assign_stmt_394_to_assign_stmt_435/MUX_434_start/req
      -- CP-element group 2: 	 assign_stmt_394_to_assign_stmt_435/call_stmt_419_update_completed_
      -- CP-element group 2: 	 assign_stmt_394_to_assign_stmt_435/call_stmt_419_Update/cca
      -- CP-element group 2: 	 assign_stmt_394_to_assign_stmt_435/call_stmt_419_Update/$exit
      -- CP-element group 2: 	 assign_stmt_394_to_assign_stmt_435/MUX_434_sample_start_
      -- 
    cca_549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_419_call_ack_1, ack => getQueueElement_CP_530_elements(2)); -- 
    req_557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_530_elements(2), ack => MUX_434_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_394_to_assign_stmt_435/MUX_434_start/ack
      -- CP-element group 3: 	 assign_stmt_394_to_assign_stmt_435/MUX_434_start/$exit
      -- CP-element group 3: 	 assign_stmt_394_to_assign_stmt_435/MUX_434_sample_completed_
      -- 
    ack_558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_434_inst_ack_0, ack => getQueueElement_CP_530_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 assign_stmt_394_to_assign_stmt_435/MUX_434_complete/$exit
      -- CP-element group 4: 	 assign_stmt_394_to_assign_stmt_435/MUX_434_complete/ack
      -- CP-element group 4: 	 assign_stmt_394_to_assign_stmt_435/$exit
      -- CP-element group 4: 	 assign_stmt_394_to_assign_stmt_435/MUX_434_update_completed_
      -- CP-element group 4: 	 $exit
      -- 
    ack_563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_434_inst_ack_1, ack => getQueueElement_CP_530_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_431_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u31_u34_403_wire : std_logic_vector(33 downto 0);
    signal NOT_u8_u8_414_wire_constant : std_logic_vector(7 downto 0);
    signal buffer_address_394 : std_logic_vector(35 downto 0);
    signal e0_423 : std_logic_vector(31 downto 0);
    signal e1_427 : std_logic_vector(31 downto 0);
    signal element_pair_419 : std_logic_vector(63 downto 0);
    signal element_pair_address_407 : std_logic_vector(35 downto 0);
    signal konst_430_wire_constant : std_logic_vector(31 downto 0);
    signal slice_399_wire : std_logic_vector(30 downto 0);
    signal type_cast_392_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_402_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_405_wire : std_logic_vector(35 downto 0);
    signal type_cast_409_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_411_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_417_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_414_wire_constant <= "11111111";
    konst_430_wire_constant <= "00000000000000000000000000000000";
    type_cast_392_wire_constant <= "000000000000000000000000000000010000";
    type_cast_402_wire_constant <= "000";
    type_cast_409_wire_constant <= "0";
    type_cast_411_wire_constant <= "1";
    type_cast_417_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    MUX_434_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_434_inst_req_0;
      MUX_434_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_434_inst_req_1;
      MUX_434_inst_ack_1<= update_ack(0);
      MUX_434_inst: SelectSplitProtocol generic map(name => "MUX_434_inst", data_width => 32, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => e1_427, y => e0_423, sel => BITSEL_u32_u1_431_wire, z => q_r_data_buffer, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through slice operator slice_399_inst
    slice_399_wire <= read_pointer_buffer(31 downto 1);
    -- flow-through slice operator slice_422_inst
    e0_423 <= element_pair_419(63 downto 32);
    -- flow-through slice operator slice_426_inst
    e1_427 <= element_pair_419(31 downto 0);
    -- interlock type_cast_405_inst
    process(CONCAT_u31_u34_403_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 33 downto 0) := CONCAT_u31_u34_403_wire(33 downto 0);
      type_cast_405_wire <= tmp_var; -- 
    end process;
    -- binary operator ADD_u36_u36_393_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, type_cast_392_wire_constant, tmp_var);
      buffer_address_394 <= tmp_var; --
    end process;
    -- binary operator ADD_u36_u36_406_inst
    process(buffer_address_394, type_cast_405_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buffer_address_394, type_cast_405_wire, tmp_var);
      element_pair_address_407 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_431_inst
    process(read_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(read_pointer_buffer, konst_430_wire_constant, tmp_var);
      BITSEL_u32_u1_431_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u31_u34_403_inst
    process(slice_399_wire) -- 
      variable tmp_var : std_logic_vector(33 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_399_wire, type_cast_402_wire_constant, tmp_var);
      CONCAT_u31_u34_403_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_419_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_419_call_req_0;
      call_stmt_419_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_419_call_req_1;
      call_stmt_419_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_409_wire_constant & type_cast_411_wire_constant & NOT_u8_u8_414_wire_constant & element_pair_address_407 & type_cast_417_wire_constant;
      element_pair_419 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getQueueElement_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity getQueuePointers is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    wp : out  std_logic_vector(31 downto 0);
    rp : out  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueuePointers;
architecture getQueuePointers_arch of getQueuePointers is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal wp_buffer :  std_logic_vector(31 downto 0);
  signal wp_update_enable: Boolean;
  signal rp_buffer :  std_logic_vector(31 downto 0);
  signal rp_update_enable: Boolean;
  signal getQueuePointers_CP_510_start: Boolean;
  signal getQueuePointers_CP_510_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_371_call_ack_0 : boolean;
  signal call_stmt_371_call_req_0 : boolean;
  signal call_stmt_371_call_ack_1 : boolean;
  signal call_stmt_371_call_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueuePointers_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueuePointers_CP_510_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueuePointers_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= wp_buffer;
  wp <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(63 downto 32) <= rp_buffer;
  rp <= out_buffer_data_out(63 downto 32);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueuePointers_CP_510_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueuePointers_CP_510_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueuePointers_CP_510_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueuePointers_CP_510: Block -- control-path 
    signal getQueuePointers_CP_510_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    getQueuePointers_CP_510_elements(0) <= getQueuePointers_CP_510_start;
    getQueuePointers_CP_510_symbol <= getQueuePointers_CP_510_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_371_to_assign_stmt_379/call_stmt_371_update_start_
      -- CP-element group 0: 	 call_stmt_371_to_assign_stmt_379/call_stmt_371_Sample/$entry
      -- CP-element group 0: 	 call_stmt_371_to_assign_stmt_379/call_stmt_371_sample_start_
      -- CP-element group 0: 	 call_stmt_371_to_assign_stmt_379/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_371_to_assign_stmt_379/call_stmt_371_Sample/crr
      -- CP-element group 0: 	 call_stmt_371_to_assign_stmt_379/call_stmt_371_Update/ccr
      -- CP-element group 0: 	 call_stmt_371_to_assign_stmt_379/call_stmt_371_Update/$entry
      -- 
    crr_523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_510_elements(0), ack => call_stmt_371_call_req_0); -- 
    ccr_528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_510_elements(0), ack => call_stmt_371_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_371_to_assign_stmt_379/call_stmt_371_sample_completed_
      -- CP-element group 1: 	 call_stmt_371_to_assign_stmt_379/call_stmt_371_Sample/cra
      -- CP-element group 1: 	 call_stmt_371_to_assign_stmt_379/call_stmt_371_Sample/$exit
      -- 
    cra_524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_371_call_ack_0, ack => getQueuePointers_CP_510_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 call_stmt_371_to_assign_stmt_379/call_stmt_371_update_completed_
      -- CP-element group 2: 	 call_stmt_371_to_assign_stmt_379/$exit
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_371_to_assign_stmt_379/call_stmt_371_Update/cca
      -- CP-element group 2: 	 call_stmt_371_to_assign_stmt_379/call_stmt_371_Update/$exit
      -- 
    cca_529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_371_call_ack_1, ack => getQueuePointers_CP_510_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_367_wire : std_logic_vector(35 downto 0);
    signal NOT_u8_u8_364_wire_constant : std_logic_vector(7 downto 0);
    signal konst_366_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_359_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_361_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_369_wire_constant : std_logic_vector(63 downto 0);
    signal wp_rp_371 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_364_wire_constant <= "11111111";
    konst_366_wire_constant <= "000000000000000000000000000000001000";
    type_cast_359_wire_constant <= "0";
    type_cast_361_wire_constant <= "1";
    type_cast_369_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- flow-through slice operator slice_374_inst
    wp_buffer <= wp_rp_371(63 downto 32);
    -- flow-through slice operator slice_378_inst
    rp_buffer <= wp_rp_371(31 downto 0);
    -- binary operator ADD_u36_u36_367_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_366_wire_constant, tmp_var);
      ADD_u36_u36_367_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_371_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_371_call_req_0;
      call_stmt_371_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_371_call_req_1;
      call_stmt_371_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_359_wire_constant & type_cast_361_wire_constant & NOT_u8_u8_364_wire_constant & ADD_u36_u36_367_wire & type_cast_369_wire_constant;
      wp_rp_371 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getQueuePointers_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity getTxPacketPointerFromServer is -- 
  generic (tag_length : integer); 
  port ( -- 
    queue_index : in  std_logic_vector(5 downto 0);
    pkt_pointer : out  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_call_data : out  std_logic_vector(36 downto 0);
    popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_return_data : in   std_logic_vector(32 downto 0);
    popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getTxPacketPointerFromServer;
architecture getTxPacketPointerFromServer_arch of getTxPacketPointerFromServer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 6)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 33)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal queue_index_buffer :  std_logic_vector(5 downto 0);
  signal queue_index_update_enable: Boolean;
  -- output port buffer signals
  signal pkt_pointer_buffer :  std_logic_vector(31 downto 0);
  signal pkt_pointer_update_enable: Boolean;
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal getTxPacketPointerFromServer_CP_2487_start: Boolean;
  signal getTxPacketPointerFromServer_CP_2487_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(67 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(31 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1274_call_ack_1 : boolean;
  signal call_stmt_1274_call_req_1 : boolean;
  signal call_stmt_1262_call_ack_1 : boolean;
  signal call_stmt_1262_call_req_1 : boolean;
  signal call_stmt_1274_call_ack_0 : boolean;
  signal call_stmt_1274_call_req_0 : boolean;
  signal call_stmt_1262_call_ack_0 : boolean;
  signal call_stmt_1262_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getTxPacketPointerFromServer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 6) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(5 downto 0) <= queue_index;
  queue_index_buffer <= in_buffer_data_out(5 downto 0);
  in_buffer_data_in(tag_length + 5 downto 6) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 5 downto 6);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 7);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= queue_index_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getTxPacketPointerFromServer_CP_2487_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getTxPacketPointerFromServer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 33) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= pkt_pointer_buffer;
  pkt_pointer <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(32 downto 32) <= status_buffer;
  status <= out_buffer_data_out(32 downto 32);
  out_buffer_data_in(tag_length + 32 downto 33) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 32 downto 33);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_2487_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  pkt_pointer_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 30) := "pkt_pointer_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_pkt_pointer_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => pkt_pointer_update_enable, clk => clk, reset => reset); --
  end block;
  status_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 25) := "status_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_status_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => status_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_2487_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_2487_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getTxPacketPointerFromServer_CP_2487: Block -- control-path 
    signal getTxPacketPointerFromServer_CP_2487_elements: BooleanArray(16 downto 0);
    -- 
  begin -- 
    getTxPacketPointerFromServer_CP_2487_elements(0) <= getTxPacketPointerFromServer_CP_2487_start;
    getTxPacketPointerFromServer_CP_2487_symbol <= getTxPacketPointerFromServer_CP_2487_elements(16);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	5 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_1252_to_stmt_1279/$entry
      -- 
    getTxPacketPointerFromServer_CP_2487_elements(1) <= getTxPacketPointerFromServer_CP_2487_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	7 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	13 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_1252_to_stmt_1279/queue_index_update_enable_out
      -- CP-element group 2: 	 assign_stmt_1252_to_stmt_1279/queue_index_update_enable
      -- 
    getTxPacketPointerFromServer_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= getTxPacketPointerFromServer_CP_2487_elements(7);
      gj_getTxPacketPointerFromServer_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2487_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	14 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	10 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_1252_to_stmt_1279/pkt_pointer_update_enable_in
      -- CP-element group 3: 	 assign_stmt_1252_to_stmt_1279/pkt_pointer_update_enable
      -- 
    getTxPacketPointerFromServer_CP_2487_elements(3) <= getTxPacketPointerFromServer_CP_2487_elements(14);
    -- CP-element group 4:  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	15 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_1252_to_stmt_1279/status_update_enable_in
      -- CP-element group 4: 	 assign_stmt_1252_to_stmt_1279/status_update_enable
      -- 
    getTxPacketPointerFromServer_CP_2487_elements(4) <= getTxPacketPointerFromServer_CP_2487_elements(15);
    -- CP-element group 5:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	1 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	7 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1262_sample_start_
      -- CP-element group 5: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1262_Sample/crr
      -- CP-element group 5: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1262_Sample/$entry
      -- 
    crr_2506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_2487_elements(5), ack => call_stmt_1262_call_req_0); -- 
    getTxPacketPointerFromServer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_2487_elements(1) & getTxPacketPointerFromServer_CP_2487_elements(7);
      gj_getTxPacketPointerFromServer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2487_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: 	11 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1262_update_start_
      -- CP-element group 6: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1262_Update/ccr
      -- CP-element group 6: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1262_Update/$entry
      -- 
    ccr_2511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_2487_elements(6), ack => call_stmt_1262_call_req_1); -- 
    getTxPacketPointerFromServer_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_2487_elements(8) & getTxPacketPointerFromServer_CP_2487_elements(11);
      gj_getTxPacketPointerFromServer_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2487_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7: marked-successors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: 	5 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1262_sample_completed_
      -- CP-element group 7: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1262_Sample/cra
      -- CP-element group 7: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1262_Sample/$exit
      -- 
    cra_2507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1262_call_ack_0, ack => getTxPacketPointerFromServer_CP_2487_elements(7)); -- 
    -- CP-element group 8:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	6 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1262_update_completed_
      -- CP-element group 8: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1262_Update/cca
      -- CP-element group 8: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1262_Update/$exit
      -- 
    cca_2512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1262_call_ack_1, ack => getTxPacketPointerFromServer_CP_2487_elements(8)); -- 
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1274_Sample/$entry
      -- CP-element group 9: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1274_sample_start_
      -- CP-element group 9: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1274_Sample/crr
      -- 
    crr_2520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_2487_elements(9), ack => call_stmt_1274_call_req_0); -- 
    getTxPacketPointerFromServer_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_2487_elements(8) & getTxPacketPointerFromServer_CP_2487_elements(11);
      gj_getTxPacketPointerFromServer_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2487_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	3 
    -- CP-element group 10: 	4 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1274_Update/ccr
      -- CP-element group 10: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1274_update_start_
      -- CP-element group 10: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1274_Update/$entry
      -- 
    ccr_2525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_2487_elements(10), ack => call_stmt_1274_call_req_1); -- 
    getTxPacketPointerFromServer_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "getTxPacketPointerFromServer_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_2487_elements(3) & getTxPacketPointerFromServer_CP_2487_elements(4) & getTxPacketPointerFromServer_CP_2487_elements(12);
      gj_getTxPacketPointerFromServer_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2487_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	6 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1274_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1274_sample_completed_
      -- CP-element group 11: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1274_Sample/cra
      -- 
    cra_2521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1274_call_ack_0, ack => getTxPacketPointerFromServer_CP_2487_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	16 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1274_Update/cca
      -- CP-element group 12: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1274_update_completed_
      -- CP-element group 12: 	 assign_stmt_1252_to_stmt_1279/call_stmt_1274_Update/$exit
      -- CP-element group 12: 	 assign_stmt_1252_to_stmt_1279/$exit
      -- 
    cca_2526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1274_call_ack_1, ack => getTxPacketPointerFromServer_CP_2487_elements(12)); -- 
    -- CP-element group 13:  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 queue_index_update_enable
      -- 
    getTxPacketPointerFromServer_CP_2487_elements(13) <= getTxPacketPointerFromServer_CP_2487_elements(2);
    -- CP-element group 14:  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	3 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 pkt_pointer_update_enable
      -- 
    -- CP-element group 15:  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	4 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 status_update_enable
      -- 
    -- CP-element group 16:  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 $exit
      -- 
    getTxPacketPointerFromServer_CP_2487_elements(16) <= getTxPacketPointerFromServer_CP_2487_elements(12);
    --  hookup: inputs to control-path 
    getTxPacketPointerFromServer_CP_2487_elements(14) <= pkt_pointer_update_enable;
    getTxPacketPointerFromServer_CP_2487_elements(15) <= status_update_enable;
    -- hookup: output from control-path 
    queue_index_update_enable <= getTxPacketPointerFromServer_CP_2487_elements(13);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u6_u6_1250_wire : std_logic_vector(5 downto 0);
    signal NOT_u4_u4_1257_wire_constant : std_logic_vector(3 downto 0);
    signal R_TX_QUEUES_REG_START_OFFSET_1249_wire_constant : std_logic_vector(5 downto 0);
    signal register_index_1252 : std_logic_vector(5 downto 0);
    signal tx_queue_pointer_32_1262 : std_logic_vector(31 downto 0);
    signal tx_queue_pointer_36_1268 : std_logic_vector(35 downto 0);
    signal type_cast_1254_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1260_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1266_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_1270_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_1257_wire_constant <= "1111";
    R_TX_QUEUES_REG_START_OFFSET_1249_wire_constant <= "001010";
    type_cast_1254_wire_constant <= "1";
    type_cast_1260_wire_constant <= "00000000000000000000000000000000";
    type_cast_1266_wire_constant <= "0000";
    type_cast_1270_wire_constant <= "1";
    -- interlock type_cast_1251_inst
    process(ADD_u6_u6_1250_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := ADD_u6_u6_1250_wire(5 downto 0);
      register_index_1252 <= tmp_var; -- 
    end process;
    -- binary operator ADD_u6_u6_1250_inst
    process(queue_index_buffer) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(queue_index_buffer, R_TX_QUEUES_REG_START_OFFSET_1249_wire_constant, tmp_var);
      ADD_u6_u6_1250_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u36_1267_inst
    process(tx_queue_pointer_32_1262) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(tx_queue_pointer_32_1262, type_cast_1266_wire_constant, tmp_var);
      tx_queue_pointer_36_1268 <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1262_call 
    AccessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1262_call_req_0;
      call_stmt_1262_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1262_call_req_1;
      call_stmt_1262_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1254_wire_constant & NOT_u4_u4_1257_wire_constant & register_index_1252 & type_cast_1260_wire_constant;
      tx_queue_pointer_32_1262 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1274_call 
    popFromQueue_call_group_1: Block -- 
      signal data_in: std_logic_vector(36 downto 0);
      signal data_out: std_logic_vector(32 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1274_call_req_0;
      call_stmt_1274_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1274_call_req_1;
      call_stmt_1274_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      popFromQueue_call_group_1_gI: SplitGuardInterface generic map(name => "popFromQueue_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1270_wire_constant & tx_queue_pointer_36_1268;
      pkt_pointer_buffer <= data_out(32 downto 1);
      status_buffer <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 37,
        owidth => 37,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => popFromQueue_call_reqs(0),
          ackR => popFromQueue_call_acks(0),
          dataR => popFromQueue_call_data(36 downto 0),
          tagR => popFromQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 33,
          owidth => 33,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => popFromQueue_return_acks(0), -- cross-over
          ackL => popFromQueue_return_reqs(0), -- cross-over
          dataL => popFromQueue_return_data(32 downto 0),
          tagL => popFromQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end getTxPacketPointerFromServer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity loadBuffer is -- 
  generic (tag_length : integer); 
  port ( -- 
    rx_buffer_pointer : in  std_logic_vector(35 downto 0);
    bad_packet_identifier : out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_data : out  std_logic_vector(51 downto 0);
    writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_data : out  std_logic_vector(35 downto 0);
    writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_data : in   std_logic_vector(35 downto 0);
    writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
    writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
    writePayloadToMem_call_data : out  std_logic_vector(71 downto 0);
    writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
    writePayloadToMem_return_data : in   std_logic_vector(16 downto 0);
    writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadBuffer;
architecture loadBuffer_arch of loadBuffer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rx_buffer_pointer_buffer :  std_logic_vector(35 downto 0);
  signal rx_buffer_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal bad_packet_identifier_buffer :  std_logic_vector(0 downto 0);
  signal bad_packet_identifier_update_enable: Boolean;
  signal loadBuffer_CP_1019_start: Boolean;
  signal loadBuffer_CP_1019_symbol: Boolean;
  -- volatile/operator module components. 
  component writeControlInformationToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buffer_pointer : in  std_logic_vector(35 downto 0);
      packet_size : in  std_logic_vector(7 downto 0);
      last_keep : in  std_logic_vector(7 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component writeEthernetHeaderToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      buf_pointer : in  std_logic_vector(35 downto 0);
      buf_position : out  std_logic_vector(35 downto 0);
      nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component writePayloadToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buf_pointer : in  std_logic_vector(35 downto 0);
      buf_pointer : in  std_logic_vector(35 downto 0);
      packet_size_32 : out  std_logic_vector(7 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      last_keep : out  std_logic_vector(7 downto 0);
      nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_710_call_req_0 : boolean;
  signal W_bad_packet_identifier_701_delayed_8_0_711_inst_ack_0 : boolean;
  signal call_stmt_701_call_ack_0 : boolean;
  signal call_stmt_701_call_ack_1 : boolean;
  signal W_rx_buffer_pointer_695_delayed_4_0_702_inst_req_1 : boolean;
  signal call_stmt_701_call_req_1 : boolean;
  signal W_bad_packet_identifier_701_delayed_8_0_711_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_695_delayed_4_0_702_inst_req_0 : boolean;
  signal call_stmt_701_call_req_0 : boolean;
  signal W_rx_buffer_pointer_702_delayed_8_0_714_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_702_delayed_8_0_714_inst_req_0 : boolean;
  signal W_rx_buffer_pointer_702_delayed_8_0_714_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_702_delayed_8_0_714_inst_ack_1 : boolean;
  signal W_rx_buffer_pointer_695_delayed_4_0_702_inst_ack_0 : boolean;
  signal call_stmt_710_call_req_1 : boolean;
  signal call_stmt_710_call_ack_0 : boolean;
  signal call_stmt_710_call_ack_1 : boolean;
  signal W_rx_buffer_pointer_695_delayed_4_0_702_inst_ack_1 : boolean;
  signal W_bad_packet_identifier_701_delayed_8_0_711_inst_ack_1 : boolean;
  signal W_bad_packet_identifier_701_delayed_8_0_711_inst_req_0 : boolean;
  signal call_stmt_721_call_req_0 : boolean;
  signal call_stmt_721_call_ack_0 : boolean;
  signal call_stmt_721_call_req_1 : boolean;
  signal call_stmt_721_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadBuffer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= rx_buffer_pointer;
  rx_buffer_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 31);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 31);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= rx_buffer_pointer_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadBuffer_CP_1019_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadBuffer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= bad_packet_identifier_buffer;
  bad_packet_identifier <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 31);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadBuffer_CP_1019_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  bad_packet_identifier_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 40) := "bad_packet_identifier_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_bad_packet_identifier_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => bad_packet_identifier_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 31,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadBuffer_CP_1019_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadBuffer_CP_1019_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadBuffer_CP_1019: Block -- control-path 
    signal loadBuffer_CP_1019_elements: BooleanArray(30 downto 0);
    -- 
  begin -- 
    loadBuffer_CP_1019_elements(0) <= loadBuffer_CP_1019_start;
    loadBuffer_CP_1019_symbol <= loadBuffer_CP_1019_elements(30);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	20 
    -- CP-element group 1: 	8 
    -- CP-element group 1: 	4 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 call_stmt_701_to_call_stmt_721/$entry
      -- 
    loadBuffer_CP_1019_elements(1) <= loadBuffer_CP_1019_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	6 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	28 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 call_stmt_701_to_call_stmt_721/rx_buffer_pointer_update_enable_out
      -- CP-element group 2: 	 call_stmt_701_to_call_stmt_721/rx_buffer_pointer_update_enable
      -- 
    loadBuffer_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1019_elements(10) & loadBuffer_CP_1019_elements(22) & loadBuffer_CP_1019_elements(6);
      gj_loadBuffer_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1019_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	29 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	13 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 call_stmt_701_to_call_stmt_721/bad_packet_identifier_update_enable
      -- CP-element group 3: 	 call_stmt_701_to_call_stmt_721/bad_packet_identifier_update_enable_in
      -- 
    loadBuffer_CP_1019_elements(3) <= loadBuffer_CP_1019_elements(29);
    -- CP-element group 4:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	6 
    -- CP-element group 4: 	27 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 call_stmt_701_to_call_stmt_721/call_stmt_701_Sample/crr
      -- CP-element group 4: 	 call_stmt_701_to_call_stmt_721/call_stmt_701_Sample/$entry
      -- CP-element group 4: 	 call_stmt_701_to_call_stmt_721/call_stmt_701_sample_start_
      -- 
    crr_1036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1019_elements(4), ack => call_stmt_701_call_req_0); -- 
    loadBuffer_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1019_elements(1) & loadBuffer_CP_1019_elements(6) & loadBuffer_CP_1019_elements(27);
      gj_loadBuffer_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1019_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	14 
    -- CP-element group 5: 	7 
    -- CP-element group 5: 	27 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_701_to_call_stmt_721/call_stmt_701_Update/$entry
      -- CP-element group 5: 	 call_stmt_701_to_call_stmt_721/call_stmt_701_Update/ccr
      -- CP-element group 5: 	 call_stmt_701_to_call_stmt_721/call_stmt_701_update_start_
      -- 
    ccr_1041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1019_elements(5), ack => call_stmt_701_call_req_1); -- 
    loadBuffer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1019_elements(14) & loadBuffer_CP_1019_elements(7) & loadBuffer_CP_1019_elements(27);
      gj_loadBuffer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1019_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: marked-successors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: 	4 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 call_stmt_701_to_call_stmt_721/call_stmt_701_Sample/cra
      -- CP-element group 6: 	 call_stmt_701_to_call_stmt_721/call_stmt_701_Sample/$exit
      -- CP-element group 6: 	 call_stmt_701_to_call_stmt_721/call_stmt_701_sample_completed_
      -- 
    cra_1037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_701_call_ack_0, ack => loadBuffer_CP_1019_elements(6)); -- 
    -- CP-element group 7:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: marked-successors 
    -- CP-element group 7: 	5 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_701_to_call_stmt_721/call_stmt_701_Update/cca
      -- CP-element group 7: 	 call_stmt_701_to_call_stmt_721/call_stmt_701_update_completed_
      -- CP-element group 7: 	 call_stmt_701_to_call_stmt_721/call_stmt_701_Update/$exit
      -- 
    cca_1042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_701_call_ack_1, ack => loadBuffer_CP_1019_elements(7)); -- 
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	10 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_701_to_call_stmt_721/assign_stmt_704_sample_start_
      -- CP-element group 8: 	 call_stmt_701_to_call_stmt_721/assign_stmt_704_Sample/$entry
      -- CP-element group 8: 	 call_stmt_701_to_call_stmt_721/assign_stmt_704_Sample/req
      -- 
    req_1050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1019_elements(8), ack => W_rx_buffer_pointer_695_delayed_4_0_702_inst_req_0); -- 
    loadBuffer_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1019_elements(1) & loadBuffer_CP_1019_elements(10);
      gj_loadBuffer_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1019_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	14 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_701_to_call_stmt_721/assign_stmt_704_update_start_
      -- CP-element group 9: 	 call_stmt_701_to_call_stmt_721/assign_stmt_704_Update/req
      -- CP-element group 9: 	 call_stmt_701_to_call_stmt_721/assign_stmt_704_Update/$entry
      -- 
    req_1055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1019_elements(9), ack => W_rx_buffer_pointer_695_delayed_4_0_702_inst_req_1); -- 
    loadBuffer_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1019_elements(11) & loadBuffer_CP_1019_elements(14);
      gj_loadBuffer_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1019_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10: marked-successors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: 	2 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_701_to_call_stmt_721/assign_stmt_704_sample_completed_
      -- CP-element group 10: 	 call_stmt_701_to_call_stmt_721/assign_stmt_704_Sample/$exit
      -- CP-element group 10: 	 call_stmt_701_to_call_stmt_721/assign_stmt_704_Sample/ack
      -- 
    ack_1051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_695_delayed_4_0_702_inst_ack_0, ack => loadBuffer_CP_1019_elements(10)); -- 
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_701_to_call_stmt_721/assign_stmt_704_update_completed_
      -- CP-element group 11: 	 call_stmt_701_to_call_stmt_721/assign_stmt_704_Update/$exit
      -- CP-element group 11: 	 call_stmt_701_to_call_stmt_721/assign_stmt_704_Update/ack
      -- 
    ack_1056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_695_delayed_4_0_702_inst_ack_1, ack => loadBuffer_CP_1019_elements(11)); -- 
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: 	7 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_701_to_call_stmt_721/call_stmt_710_sample_start_
      -- CP-element group 12: 	 call_stmt_701_to_call_stmt_721/call_stmt_710_Sample/crr
      -- CP-element group 12: 	 call_stmt_701_to_call_stmt_721/call_stmt_710_Sample/$entry
      -- 
    crr_1064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1019_elements(12), ack => call_stmt_710_call_req_0); -- 
    loadBuffer_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1019_elements(11) & loadBuffer_CP_1019_elements(7) & loadBuffer_CP_1019_elements(14);
      gj_loadBuffer_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1019_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	3 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: 	18 
    -- CP-element group 13: 	26 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_701_to_call_stmt_721/call_stmt_710_Update/$entry
      -- CP-element group 13: 	 call_stmt_701_to_call_stmt_721/call_stmt_710_update_start_
      -- CP-element group 13: 	 call_stmt_701_to_call_stmt_721/call_stmt_710_Update/ccr
      -- 
    ccr_1069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1019_elements(13), ack => call_stmt_710_call_req_1); -- 
    loadBuffer_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= loadBuffer_CP_1019_elements(3) & loadBuffer_CP_1019_elements(15) & loadBuffer_CP_1019_elements(18) & loadBuffer_CP_1019_elements(26);
      gj_loadBuffer_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1019_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: 	9 
    -- CP-element group 14: 	5 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 call_stmt_701_to_call_stmt_721/call_stmt_710_sample_completed_
      -- CP-element group 14: 	 call_stmt_701_to_call_stmt_721/call_stmt_710_Sample/$exit
      -- CP-element group 14: 	 call_stmt_701_to_call_stmt_721/call_stmt_710_Sample/cra
      -- 
    cra_1065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_710_call_ack_0, ack => loadBuffer_CP_1019_elements(14)); -- 
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	24 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	13 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 call_stmt_701_to_call_stmt_721/call_stmt_710_Update/$exit
      -- CP-element group 15: 	 call_stmt_701_to_call_stmt_721/call_stmt_710_update_completed_
      -- CP-element group 15: 	 call_stmt_701_to_call_stmt_721/call_stmt_710_Update/cca
      -- 
    cca_1070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_710_call_ack_1, ack => loadBuffer_CP_1019_elements(15)); -- 
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	18 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 call_stmt_701_to_call_stmt_721/assign_stmt_713_Sample/$entry
      -- CP-element group 16: 	 call_stmt_701_to_call_stmt_721/assign_stmt_713_sample_start_
      -- CP-element group 16: 	 call_stmt_701_to_call_stmt_721/assign_stmt_713_Sample/req
      -- 
    req_1078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1019_elements(16), ack => W_bad_packet_identifier_701_delayed_8_0_711_inst_req_0); -- 
    loadBuffer_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1019_elements(15) & loadBuffer_CP_1019_elements(18);
      gj_loadBuffer_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1019_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: 	26 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 call_stmt_701_to_call_stmt_721/assign_stmt_713_Update/$entry
      -- CP-element group 17: 	 call_stmt_701_to_call_stmt_721/assign_stmt_713_Update/req
      -- CP-element group 17: 	 call_stmt_701_to_call_stmt_721/assign_stmt_713_update_start_
      -- 
    req_1083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1019_elements(17), ack => W_bad_packet_identifier_701_delayed_8_0_711_inst_req_1); -- 
    loadBuffer_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1019_elements(19) & loadBuffer_CP_1019_elements(26);
      gj_loadBuffer_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1019_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	13 
    -- CP-element group 18: 	16 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 call_stmt_701_to_call_stmt_721/assign_stmt_713_Sample/ack
      -- CP-element group 18: 	 call_stmt_701_to_call_stmt_721/assign_stmt_713_Sample/$exit
      -- CP-element group 18: 	 call_stmt_701_to_call_stmt_721/assign_stmt_713_sample_completed_
      -- 
    ack_1079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bad_packet_identifier_701_delayed_8_0_711_inst_ack_0, ack => loadBuffer_CP_1019_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	24 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	17 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 call_stmt_701_to_call_stmt_721/assign_stmt_713_Update/$exit
      -- CP-element group 19: 	 call_stmt_701_to_call_stmt_721/assign_stmt_713_update_completed_
      -- CP-element group 19: 	 call_stmt_701_to_call_stmt_721/assign_stmt_713_Update/ack
      -- 
    ack_1084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bad_packet_identifier_701_delayed_8_0_711_inst_ack_1, ack => loadBuffer_CP_1019_elements(19)); -- 
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	1 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	22 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 call_stmt_701_to_call_stmt_721/assign_stmt_716_sample_start_
      -- CP-element group 20: 	 call_stmt_701_to_call_stmt_721/assign_stmt_716_Sample/req
      -- CP-element group 20: 	 call_stmt_701_to_call_stmt_721/assign_stmt_716_Sample/$entry
      -- 
    req_1092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1019_elements(20), ack => W_rx_buffer_pointer_702_delayed_8_0_714_inst_req_0); -- 
    loadBuffer_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1019_elements(1) & loadBuffer_CP_1019_elements(22);
      gj_loadBuffer_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1019_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: 	26 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 call_stmt_701_to_call_stmt_721/assign_stmt_716_update_start_
      -- CP-element group 21: 	 call_stmt_701_to_call_stmt_721/assign_stmt_716_Update/$entry
      -- CP-element group 21: 	 call_stmt_701_to_call_stmt_721/assign_stmt_716_Update/req
      -- 
    req_1097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1019_elements(21), ack => W_rx_buffer_pointer_702_delayed_8_0_714_inst_req_1); -- 
    loadBuffer_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1019_elements(23) & loadBuffer_CP_1019_elements(26);
      gj_loadBuffer_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1019_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: 	2 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 call_stmt_701_to_call_stmt_721/assign_stmt_716_sample_completed_
      -- CP-element group 22: 	 call_stmt_701_to_call_stmt_721/assign_stmt_716_Sample/ack
      -- CP-element group 22: 	 call_stmt_701_to_call_stmt_721/assign_stmt_716_Sample/$exit
      -- 
    ack_1093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_702_delayed_8_0_714_inst_ack_0, ack => loadBuffer_CP_1019_elements(22)); -- 
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	21 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 call_stmt_701_to_call_stmt_721/assign_stmt_716_update_completed_
      -- CP-element group 23: 	 call_stmt_701_to_call_stmt_721/assign_stmt_716_Update/$exit
      -- CP-element group 23: 	 call_stmt_701_to_call_stmt_721/assign_stmt_716_Update/ack
      -- 
    ack_1098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_702_delayed_8_0_714_inst_ack_1, ack => loadBuffer_CP_1019_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	15 
    -- CP-element group 24: 	19 
    -- CP-element group 24: 	23 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 call_stmt_701_to_call_stmt_721/call_stmt_721_sample_start_
      -- CP-element group 24: 	 call_stmt_701_to_call_stmt_721/call_stmt_721_Sample/$entry
      -- CP-element group 24: 	 call_stmt_701_to_call_stmt_721/call_stmt_721_Sample/crr
      -- 
    crr_1106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1019_elements(24), ack => call_stmt_721_call_req_0); -- 
    loadBuffer_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= loadBuffer_CP_1019_elements(15) & loadBuffer_CP_1019_elements(19) & loadBuffer_CP_1019_elements(23) & loadBuffer_CP_1019_elements(26);
      gj_loadBuffer_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1019_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	27 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 call_stmt_701_to_call_stmt_721/call_stmt_721_update_start_
      -- CP-element group 25: 	 call_stmt_701_to_call_stmt_721/call_stmt_721_Update/$entry
      -- CP-element group 25: 	 call_stmt_701_to_call_stmt_721/call_stmt_721_Update/ccr
      -- 
    ccr_1111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1019_elements(25), ack => call_stmt_721_call_req_1); -- 
    loadBuffer_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= loadBuffer_CP_1019_elements(27);
      gj_loadBuffer_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1019_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	13 
    -- CP-element group 26: 	17 
    -- CP-element group 26: 	21 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 call_stmt_701_to_call_stmt_721/call_stmt_721_sample_completed_
      -- CP-element group 26: 	 call_stmt_701_to_call_stmt_721/call_stmt_721_Sample/$exit
      -- CP-element group 26: 	 call_stmt_701_to_call_stmt_721/call_stmt_721_Sample/cra
      -- 
    cra_1107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_721_call_ack_0, ack => loadBuffer_CP_1019_elements(26)); -- 
    -- CP-element group 27:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	30 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: 	4 
    -- CP-element group 27: 	5 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 call_stmt_701_to_call_stmt_721/$exit
      -- CP-element group 27: 	 call_stmt_701_to_call_stmt_721/call_stmt_721_update_completed_
      -- CP-element group 27: 	 call_stmt_701_to_call_stmt_721/call_stmt_721_Update/$exit
      -- CP-element group 27: 	 call_stmt_701_to_call_stmt_721/call_stmt_721_Update/cca
      -- 
    cca_1112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_721_call_ack_1, ack => loadBuffer_CP_1019_elements(27)); -- 
    -- CP-element group 28:  place  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 rx_buffer_pointer_update_enable
      -- 
    loadBuffer_CP_1019_elements(28) <= loadBuffer_CP_1019_elements(2);
    -- CP-element group 29:  place  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	3 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 bad_packet_identifier_update_enable
      -- 
    -- CP-element group 30:  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 $exit
      -- 
    loadBuffer_CP_1019_elements(30) <= loadBuffer_CP_1019_elements(27);
    --  hookup: inputs to control-path 
    loadBuffer_CP_1019_elements(29) <= bad_packet_identifier_update_enable;
    -- hookup: output from control-path 
    rx_buffer_pointer_update_enable <= loadBuffer_CP_1019_elements(28);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal bad_packet_identifier_701_delayed_8_0_713 : std_logic_vector(0 downto 0);
    signal last_keep_710 : std_logic_vector(7 downto 0);
    signal new_buf_pointer_701 : std_logic_vector(35 downto 0);
    signal packet_size_710 : std_logic_vector(7 downto 0);
    signal rx_buffer_pointer_695_delayed_4_0_704 : std_logic_vector(35 downto 0);
    signal rx_buffer_pointer_702_delayed_8_0_716 : std_logic_vector(35 downto 0);
    -- 
  begin -- 
    W_bad_packet_identifier_701_delayed_8_0_711_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_bad_packet_identifier_701_delayed_8_0_711_inst_req_0;
      W_bad_packet_identifier_701_delayed_8_0_711_inst_ack_0<= wack(0);
      rreq(0) <= W_bad_packet_identifier_701_delayed_8_0_711_inst_req_1;
      W_bad_packet_identifier_701_delayed_8_0_711_inst_ack_1<= rack(0);
      W_bad_packet_identifier_701_delayed_8_0_711_inst : InterlockBuffer generic map ( -- 
        name => "W_bad_packet_identifier_701_delayed_8_0_711_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => bad_packet_identifier_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => bad_packet_identifier_701_delayed_8_0_713,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_695_delayed_4_0_702_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_695_delayed_4_0_702_inst_req_0;
      W_rx_buffer_pointer_695_delayed_4_0_702_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_695_delayed_4_0_702_inst_req_1;
      W_rx_buffer_pointer_695_delayed_4_0_702_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_695_delayed_4_0_702_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_695_delayed_4_0_702_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_695_delayed_4_0_704,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_702_delayed_8_0_714_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_702_delayed_8_0_714_inst_req_0;
      W_rx_buffer_pointer_702_delayed_8_0_714_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_702_delayed_8_0_714_inst_req_1;
      W_rx_buffer_pointer_702_delayed_8_0_714_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_702_delayed_8_0_714_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_702_delayed_8_0_714_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_702_delayed_8_0_716,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- shared call operator group (0) : call_stmt_701_call 
    writeEthernetHeaderToMem_call_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_701_call_req_0;
      call_stmt_701_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_701_call_req_1;
      call_stmt_701_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeEthernetHeaderToMem_call_group_0_gI: SplitGuardInterface generic map(name => "writeEthernetHeaderToMem_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_buffer;
      new_buf_pointer_701 <= data_out(35 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeEthernetHeaderToMem_call_reqs(0),
          ackR => writeEthernetHeaderToMem_call_acks(0),
          dataR => writeEthernetHeaderToMem_call_data(35 downto 0),
          tagR => writeEthernetHeaderToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 36,
          owidth => 36,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => writeEthernetHeaderToMem_return_acks(0), -- cross-over
          ackL => writeEthernetHeaderToMem_return_reqs(0), -- cross-over
          dataL => writeEthernetHeaderToMem_return_data(35 downto 0),
          tagL => writeEthernetHeaderToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_710_call 
    writePayloadToMem_call_group_1: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(16 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_710_call_req_0;
      call_stmt_710_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_710_call_req_1;
      call_stmt_710_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writePayloadToMem_call_group_1_gI: SplitGuardInterface generic map(name => "writePayloadToMem_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_695_delayed_4_0_704 & new_buf_pointer_701;
      packet_size_710 <= data_out(16 downto 9);
      bad_packet_identifier_buffer <= data_out(8 downto 8);
      last_keep_710 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writePayloadToMem_call_reqs(0),
          ackR => writePayloadToMem_call_acks(0),
          dataR => writePayloadToMem_call_data(71 downto 0),
          tagR => writePayloadToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 17,
          owidth => 17,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => writePayloadToMem_return_acks(0), -- cross-over
          ackL => writePayloadToMem_return_reqs(0), -- cross-over
          dataL => writePayloadToMem_return_data(16 downto 0),
          tagL => writePayloadToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_721_call 
    writeControlInformationToMem_call_group_2: Block -- 
      signal data_in: std_logic_vector(51 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_721_call_req_0;
      call_stmt_721_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_721_call_req_1;
      call_stmt_721_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not bad_packet_identifier_701_delayed_8_0_713(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeControlInformationToMem_call_group_2_gI: SplitGuardInterface generic map(name => "writeControlInformationToMem_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_702_delayed_8_0_716 & packet_size_710 & last_keep_710;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 52,
        owidth => 52,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeControlInformationToMem_call_reqs(0),
          ackR => writeControlInformationToMem_call_acks(0),
          dataR => writeControlInformationToMem_call_data(51 downto 0),
          tagR => writeControlInformationToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => writeControlInformationToMem_return_acks(0), -- cross-over
          ackL => writeControlInformationToMem_return_reqs(0), -- cross-over
          tagL => writeControlInformationToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end loadBuffer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity nextLSTATE_Volatile is -- 
  port ( -- 
    RX : in  std_logic_vector(72 downto 0);
    LSTATE : in  std_logic_vector(1 downto 0);
    nLSTATE : out  std_logic_vector(1 downto 0)-- 
  );
  -- 
end entity nextLSTATE_Volatile;
architecture nextLSTATE_Volatile_arch of nextLSTATE_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(75-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal RX_buffer :  std_logic_vector(72 downto 0);
  signal LSTATE_buffer :  std_logic_vector(1 downto 0);
  -- output port buffer signals
  signal nLSTATE_buffer :  std_logic_vector(1 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  RX_buffer <= RX;
  LSTATE_buffer <= LSTATE;
  -- output handling  -------------------------------------------------------
  nLSTATE <= nLSTATE_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_1316_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1324_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1300_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1306_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1313_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1322_wire : std_logic_vector(0 downto 0);
    signal MUX_1303_wire : std_logic_vector(1 downto 0);
    signal MUX_1309_wire : std_logic_vector(1 downto 0);
    signal MUX_1319_wire : std_logic_vector(1 downto 0);
    signal MUX_1327_wire : std_logic_vector(1 downto 0);
    signal NOT_u1_u1_1315_wire : std_logic_vector(0 downto 0);
    signal OR_u2_u2_1310_wire : std_logic_vector(1 downto 0);
    signal OR_u2_u2_1328_wire : std_logic_vector(1 downto 0);
    signal R_S0_1299_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_1325_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_1301_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_1305_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1307_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1312_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1317_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1321_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1294_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1302_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1308_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1318_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1326_wire_constant : std_logic_vector(1 downto 0);
    signal last_word_1296 : std_logic_vector(0 downto 0);
    signal tlast_1291 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_S0_1299_wire_constant <= "00";
    R_S0_1325_wire_constant <= "00";
    R_S1_1301_wire_constant <= "01";
    R_S1_1305_wire_constant <= "01";
    R_S2_1307_wire_constant <= "10";
    R_S2_1312_wire_constant <= "10";
    R_S2_1317_wire_constant <= "10";
    R_S2_1321_wire_constant <= "10";
    konst_1294_wire_constant <= "1";
    konst_1302_wire_constant <= "00";
    konst_1308_wire_constant <= "00";
    konst_1318_wire_constant <= "00";
    konst_1326_wire_constant <= "00";
    -- flow-through select operator MUX_1303_inst
    MUX_1303_wire <= R_S1_1301_wire_constant when (EQ_u2_u1_1300_wire(0) /=  '0') else konst_1302_wire_constant;
    -- flow-through select operator MUX_1309_inst
    MUX_1309_wire <= R_S2_1307_wire_constant when (EQ_u2_u1_1306_wire(0) /=  '0') else konst_1308_wire_constant;
    -- flow-through select operator MUX_1319_inst
    MUX_1319_wire <= R_S2_1317_wire_constant when (AND_u1_u1_1316_wire(0) /=  '0') else konst_1318_wire_constant;
    -- flow-through select operator MUX_1327_inst
    MUX_1327_wire <= R_S0_1325_wire_constant when (AND_u1_u1_1324_wire(0) /=  '0') else konst_1326_wire_constant;
    -- flow-through slice operator slice_1290_inst
    tlast_1291 <= RX_buffer(72 downto 72);
    -- binary operator AND_u1_u1_1316_inst
    process(EQ_u2_u1_1313_wire, NOT_u1_u1_1315_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_1313_wire, NOT_u1_u1_1315_wire, tmp_var);
      AND_u1_u1_1316_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1324_inst
    process(EQ_u2_u1_1322_wire, last_word_1296) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_1322_wire, last_word_1296, tmp_var);
      AND_u1_u1_1324_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1295_inst
    process(tlast_1291) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(tlast_1291, konst_1294_wire_constant, tmp_var);
      last_word_1296 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1300_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S0_1299_wire_constant, tmp_var);
      EQ_u2_u1_1300_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1306_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S1_1305_wire_constant, tmp_var);
      EQ_u2_u1_1306_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1313_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S2_1312_wire_constant, tmp_var);
      EQ_u2_u1_1313_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1322_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S2_1321_wire_constant, tmp_var);
      EQ_u2_u1_1322_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1315_inst
    process(last_word_1296) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", last_word_1296, tmp_var);
      NOT_u1_u1_1315_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u2_u2_1310_inst
    process(MUX_1303_wire, MUX_1309_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1303_wire, MUX_1309_wire, tmp_var);
      OR_u2_u2_1310_wire <= tmp_var; --
    end process;
    -- binary operator OR_u2_u2_1328_inst
    process(MUX_1319_wire, MUX_1327_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1319_wire, MUX_1327_wire, tmp_var);
      OR_u2_u2_1328_wire <= tmp_var; --
    end process;
    -- binary operator OR_u2_u2_1329_inst
    process(OR_u2_u2_1310_wire, OR_u2_u2_1328_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u2_u2_1310_wire, OR_u2_u2_1328_wire, tmp_var);
      nLSTATE_buffer <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end nextLSTATE_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity nicRxFromMacDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    mac_to_nic_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_read_data : in   std_logic_vector(72 downto 0);
    CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    nic_rx_to_packet_pipe_write_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_write_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_write_data : out  std_logic_vector(72 downto 0);
    nic_rx_to_header_pipe_write_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_write_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_write_data : out  std_logic_vector(72 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity nicRxFromMacDaemon;
architecture nicRxFromMacDaemon_arch of nicRxFromMacDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal nicRxFromMacDaemon_CP_2536_start: Boolean;
  signal nicRxFromMacDaemon_CP_2536_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component nextLSTATE_Volatile is -- 
    port ( -- 
      RX : in  std_logic_vector(72 downto 0);
      LSTATE : in  std_logic_vector(1 downto 0);
      nLSTATE : out  std_logic_vector(1 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal do_while_stmt_1364_branch_ack_0 : boolean;
  signal WPIPE_nic_rx_to_packet_1402_inst_ack_0 : boolean;
  signal WPIPE_nic_rx_to_packet_1402_inst_req_0 : boolean;
  signal WPIPE_nic_rx_to_packet_1402_inst_req_1 : boolean;
  signal do_while_stmt_1364_branch_ack_1 : boolean;
  signal WPIPE_nic_rx_to_packet_1402_inst_ack_1 : boolean;
  signal call_stmt_1345_call_req_0 : boolean;
  signal call_stmt_1345_call_ack_0 : boolean;
  signal call_stmt_1345_call_req_1 : boolean;
  signal call_stmt_1345_call_ack_1 : boolean;
  signal if_stmt_1346_branch_req_0 : boolean;
  signal if_stmt_1346_branch_ack_1 : boolean;
  signal if_stmt_1346_branch_ack_0 : boolean;
  signal call_stmt_1363_call_req_0 : boolean;
  signal call_stmt_1363_call_ack_0 : boolean;
  signal call_stmt_1363_call_req_1 : boolean;
  signal call_stmt_1363_call_ack_1 : boolean;
  signal do_while_stmt_1364_branch_req_0 : boolean;
  signal phi_stmt_1366_req_0 : boolean;
  signal phi_stmt_1366_req_1 : boolean;
  signal phi_stmt_1366_ack_0 : boolean;
  signal nLSTATE_1380_1368_buf_req_0 : boolean;
  signal nLSTATE_1380_1368_buf_ack_0 : boolean;
  signal nLSTATE_1380_1368_buf_req_1 : boolean;
  signal nLSTATE_1380_1368_buf_ack_1 : boolean;
  signal RPIPE_mac_to_nic_data_1372_inst_req_0 : boolean;
  signal RPIPE_mac_to_nic_data_1372_inst_ack_0 : boolean;
  signal RPIPE_mac_to_nic_data_1372_inst_req_1 : boolean;
  signal RPIPE_mac_to_nic_data_1372_inst_ack_1 : boolean;
  signal MUX_1400_inst_req_0 : boolean;
  signal MUX_1400_inst_ack_0 : boolean;
  signal MUX_1400_inst_req_1 : boolean;
  signal MUX_1400_inst_ack_1 : boolean;
  signal WPIPE_nic_rx_to_header_1391_inst_req_0 : boolean;
  signal WPIPE_nic_rx_to_header_1391_inst_ack_0 : boolean;
  signal WPIPE_nic_rx_to_header_1391_inst_req_1 : boolean;
  signal WPIPE_nic_rx_to_header_1391_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "nicRxFromMacDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  nicRxFromMacDaemon_CP_2536_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "nicRxFromMacDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_2536_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_2536_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_2536_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  nicRxFromMacDaemon_CP_2536: Block -- control-path 
    signal nicRxFromMacDaemon_CP_2536_elements: BooleanArray(59 downto 0);
    -- 
  begin -- 
    nicRxFromMacDaemon_CP_2536_elements(0) <= nicRxFromMacDaemon_CP_2536_start;
    nicRxFromMacDaemon_CP_2536_symbol <= nicRxFromMacDaemon_CP_2536_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	59 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 branch_block_stmt_1333/merge_stmt_1335__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_1333/merge_stmt_1335__entry___PhiReq/$exit
      -- CP-element group 0: 	 branch_block_stmt_1333/merge_stmt_1335_dead_link/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1333/$entry
      -- CP-element group 0: 	 branch_block_stmt_1333/branch_block_stmt_1333__entry__
      -- CP-element group 0: 	 branch_block_stmt_1333/merge_stmt_1335__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1333/$exit
      -- CP-element group 1: 	 branch_block_stmt_1333/branch_block_stmt_1333__exit__
      -- 
    nicRxFromMacDaemon_CP_2536_elements(1) <= false; 
    -- CP-element group 2:  transition  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	58 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	59 
    -- CP-element group 2:  members (4) 
      -- CP-element group 2: 	 branch_block_stmt_1333/disable_loopback_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_1333/disable_loopback_PhiReq/$exit
      -- CP-element group 2: 	 branch_block_stmt_1333/do_while_stmt_1364__exit__
      -- CP-element group 2: 	 branch_block_stmt_1333/disable_loopback
      -- 
    nicRxFromMacDaemon_CP_2536_elements(2) <= nicRxFromMacDaemon_CP_2536_elements(58);
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	59 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1333/call_stmt_1345/call_stmt_1345_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1333/call_stmt_1345/call_stmt_1345_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1333/call_stmt_1345/call_stmt_1345_Sample/cra
      -- 
    cra_2566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1345_call_ack_0, ack => nicRxFromMacDaemon_CP_2536_elements(3)); -- 
    -- CP-element group 4:  branch  transition  place  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	59 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (49) 
      -- CP-element group 4: 	 branch_block_stmt_1333/call_stmt_1345__exit__
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346__entry__
      -- CP-element group 4: 	 branch_block_stmt_1333/call_stmt_1345/$exit
      -- CP-element group 4: 	 branch_block_stmt_1333/call_stmt_1345/call_stmt_1345_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1333/call_stmt_1345/call_stmt_1345_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1333/call_stmt_1345/call_stmt_1345_Update/cca
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_dead_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/$entry
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/$exit
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/$entry
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/$exit
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/$entry
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/$exit
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/BITSEL_u32_u1_1349_inputs/$entry
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/BITSEL_u32_u1_1349_inputs/$exit
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/BITSEL_u32_u1_1349_inputs/RPIPE_CONTROL_REGISTER_1347/$entry
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/BITSEL_u32_u1_1349_inputs/RPIPE_CONTROL_REGISTER_1347/$exit
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/BITSEL_u32_u1_1349_inputs/RPIPE_CONTROL_REGISTER_1347/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/BITSEL_u32_u1_1349_inputs/RPIPE_CONTROL_REGISTER_1347/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/BITSEL_u32_u1_1349_inputs/RPIPE_CONTROL_REGISTER_1347/Sample/req
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/BITSEL_u32_u1_1349_inputs/RPIPE_CONTROL_REGISTER_1347/Sample/ack
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/BITSEL_u32_u1_1349_inputs/RPIPE_CONTROL_REGISTER_1347/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/BITSEL_u32_u1_1349_inputs/RPIPE_CONTROL_REGISTER_1347/Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/BITSEL_u32_u1_1349_inputs/RPIPE_CONTROL_REGISTER_1347/Update/req
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/BITSEL_u32_u1_1349_inputs/RPIPE_CONTROL_REGISTER_1347/Update/ack
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/SplitProtocol/$exit
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/SplitProtocol/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/SplitProtocol/Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/SplitProtocol/Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/BITSEL_u32_u1_1349/SplitProtocol/Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/SplitProtocol/$exit
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/SplitProtocol/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/SplitProtocol/Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/SplitProtocol/Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/NOT_u1_u1_1350/SplitProtocol/Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_eval_test/branch_req
      -- CP-element group 4: 	 branch_block_stmt_1333/NOT_u1_u1_1350_place
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_if_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_1333/if_stmt_1346_else_link/$entry
      -- 
    cca_2571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1345_call_ack_1, ack => nicRxFromMacDaemon_CP_2536_elements(4)); -- 
    branch_req_2627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2536_elements(4), ack => if_stmt_1346_branch_req_0); -- 
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	59 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1333/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_1333/not_enabled_yet_loopback_PhiReq/$exit
      -- CP-element group 5: 	 branch_block_stmt_1333/if_stmt_1346_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_1333/if_stmt_1346_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_1333/not_enabled_yet_loopback
      -- 
    if_choice_transition_2632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1346_branch_ack_1, ack => nicRxFromMacDaemon_CP_2536_elements(5)); -- 
    -- CP-element group 6:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_1333/if_stmt_1346__exit__
      -- CP-element group 6: 	 branch_block_stmt_1333/call_stmt_1363__entry__
      -- CP-element group 6: 	 branch_block_stmt_1333/if_stmt_1346_else_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_1333/if_stmt_1346_else_link/else_choice_transition
      -- CP-element group 6: 	 branch_block_stmt_1333/call_stmt_1363/$entry
      -- CP-element group 6: 	 branch_block_stmt_1333/call_stmt_1363/call_stmt_1363_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1333/call_stmt_1363/call_stmt_1363_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1333/call_stmt_1363/call_stmt_1363_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1333/call_stmt_1363/call_stmt_1363_Sample/crr
      -- CP-element group 6: 	 branch_block_stmt_1333/call_stmt_1363/call_stmt_1363_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1333/call_stmt_1363/call_stmt_1363_Update/ccr
      -- 
    else_choice_transition_2636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1346_branch_ack_0, ack => nicRxFromMacDaemon_CP_2536_elements(6)); -- 
    crr_2648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2536_elements(6), ack => call_stmt_1363_call_req_0); -- 
    ccr_2653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2536_elements(6), ack => call_stmt_1363_call_req_1); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1333/call_stmt_1363/call_stmt_1363_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1333/call_stmt_1363/call_stmt_1363_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1333/call_stmt_1363/call_stmt_1363_Sample/cra
      -- 
    cra_2649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1363_call_ack_0, ack => nicRxFromMacDaemon_CP_2536_elements(7)); -- 
    -- CP-element group 8:  transition  place  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1333/call_stmt_1363__exit__
      -- CP-element group 8: 	 branch_block_stmt_1333/do_while_stmt_1364__entry__
      -- CP-element group 8: 	 branch_block_stmt_1333/call_stmt_1363/$exit
      -- CP-element group 8: 	 branch_block_stmt_1333/call_stmt_1363/call_stmt_1363_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1333/call_stmt_1363/call_stmt_1363_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1333/call_stmt_1363/call_stmt_1363_Update/cca
      -- 
    cca_2654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1363_call_ack_1, ack => nicRxFromMacDaemon_CP_2536_elements(8)); -- 
    -- CP-element group 9:  transition  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	15 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1333/do_while_stmt_1364/$entry
      -- CP-element group 9: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364__entry__
      -- 
    nicRxFromMacDaemon_CP_2536_elements(9) <= nicRxFromMacDaemon_CP_2536_elements(8);
    -- CP-element group 10:  merge  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	58 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364__exit__
      -- 
    -- Element group nicRxFromMacDaemon_CP_2536_elements(10) is bound as output of CP function.
    -- CP-element group 11:  merge  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1333/do_while_stmt_1364/loop_back
      -- 
    -- Element group nicRxFromMacDaemon_CP_2536_elements(11) is bound as output of CP function.
    -- CP-element group 12:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	56 
    -- CP-element group 12: 	57 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1333/do_while_stmt_1364/loop_taken/$entry
      -- CP-element group 12: 	 branch_block_stmt_1333/do_while_stmt_1364/loop_exit/$entry
      -- CP-element group 12: 	 branch_block_stmt_1333/do_while_stmt_1364/condition_done
      -- 
    nicRxFromMacDaemon_CP_2536_elements(12) <= nicRxFromMacDaemon_CP_2536_elements(17);
    -- CP-element group 13:  branch  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	55 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1333/do_while_stmt_1364/loop_body_done
      -- 
    nicRxFromMacDaemon_CP_2536_elements(13) <= nicRxFromMacDaemon_CP_2536_elements(55);
    -- CP-element group 14:  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	26 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/back_edge_to_loop_body
      -- 
    nicRxFromMacDaemon_CP_2536_elements(14) <= nicRxFromMacDaemon_CP_2536_elements(11);
    -- CP-element group 15:  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	28 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/first_time_through_loop_body
      -- 
    nicRxFromMacDaemon_CP_2536_elements(15) <= nicRxFromMacDaemon_CP_2536_elements(9);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	39 
    -- CP-element group 16: 	18 
    -- CP-element group 16: 	22 
    -- CP-element group 16: 	23 
    -- CP-element group 16: 	54 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/$entry
      -- CP-element group 16: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/loop_body_start
      -- CP-element group 16: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1370_sample_start_
      -- 
    -- Element group nicRxFromMacDaemon_CP_2536_elements(16) is bound as output of CP function.
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	21 
    -- CP-element group 17: 	54 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/condition_evaluated
      -- 
    condition_evaluated_2669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2536_elements(17), ack => do_while_stmt_1364_branch_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2536_elements(21) & nicRxFromMacDaemon_CP_2536_elements(54);
      gj_nicRxFromMacDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2536_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: 	22 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	21 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	40 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/aggregated_phi_sample_req
      -- CP-element group 18: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1366_sample_start__ps
      -- 
    nicRxFromMacDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2536_elements(16) & nicRxFromMacDaemon_CP_2536_elements(22) & nicRxFromMacDaemon_CP_2536_elements(21);
      gj_nicRxFromMacDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2536_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	42 
    -- CP-element group 19: 	24 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	55 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/aggregated_phi_sample_ack
      -- CP-element group 19: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1366_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1370_sample_completed_
      -- 
    nicRxFromMacDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2536_elements(42) & nicRxFromMacDaemon_CP_2536_elements(24);
      gj_nicRxFromMacDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2536_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	39 
    -- CP-element group 20: 	23 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	41 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/aggregated_phi_update_req
      -- CP-element group 20: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1366_update_start__ps
      -- 
    nicRxFromMacDaemon_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2536_elements(39) & nicRxFromMacDaemon_CP_2536_elements(23);
      gj_nicRxFromMacDaemon_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2536_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	43 
    -- CP-element group 21: 	25 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	17 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	18 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/aggregated_phi_update_ack
      -- 
    nicRxFromMacDaemon_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2536_elements(43) & nicRxFromMacDaemon_CP_2536_elements(25);
      gj_nicRxFromMacDaemon_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2536_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	16 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	18 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1366_sample_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2536_elements(16) & nicRxFromMacDaemon_CP_2536_elements(19);
      gj_nicRxFromMacDaemon_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2536_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	16 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	46 
    -- CP-element group 23: 	25 
    -- CP-element group 23: 	49 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1366_update_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2536_elements(16) & nicRxFromMacDaemon_CP_2536_elements(46) & nicRxFromMacDaemon_CP_2536_elements(25) & nicRxFromMacDaemon_CP_2536_elements(49);
      gj_nicRxFromMacDaemon_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2536_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	19 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1366_sample_completed__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_2536_elements(24) is bound as output of CP function.
    -- CP-element group 25:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	44 
    -- CP-element group 25: 	21 
    -- CP-element group 25: 	48 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1366_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1366_update_completed__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_2536_elements(25) is bound as output of CP function.
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	14 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1366_loopback_trigger
      -- 
    nicRxFromMacDaemon_CP_2536_elements(26) <= nicRxFromMacDaemon_CP_2536_elements(14);
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1366_loopback_sample_req
      -- CP-element group 27: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1366_loopback_sample_req_ps
      -- 
    phi_stmt_1366_loopback_sample_req_2684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1366_loopback_sample_req_2684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2536_elements(27), ack => phi_stmt_1366_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_2536_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	15 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1366_entry_trigger
      -- 
    nicRxFromMacDaemon_CP_2536_elements(28) <= nicRxFromMacDaemon_CP_2536_elements(15);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1366_entry_sample_req
      -- CP-element group 29: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1366_entry_sample_req_ps
      -- 
    phi_stmt_1366_entry_sample_req_2687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1366_entry_sample_req_2687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2536_elements(29), ack => phi_stmt_1366_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_2536_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1366_phi_mux_ack
      -- CP-element group 30: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1366_phi_mux_ack_ps
      -- 
    phi_stmt_1366_phi_mux_ack_2690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1366_ack_0, ack => nicRxFromMacDaemon_CP_2536_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_nLSTATE_1368_sample_start__ps
      -- CP-element group 31: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_nLSTATE_1368_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_nLSTATE_1368_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_nLSTATE_1368_Sample/req
      -- 
    req_2703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2536_elements(31), ack => nLSTATE_1380_1368_buf_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_2536_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_nLSTATE_1368_update_start__ps
      -- CP-element group 32: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_nLSTATE_1368_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_nLSTATE_1368_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_nLSTATE_1368_Update/req
      -- 
    req_2708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2536_elements(32), ack => nLSTATE_1380_1368_buf_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_2536_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_nLSTATE_1368_sample_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_nLSTATE_1368_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_nLSTATE_1368_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_nLSTATE_1368_Sample/ack
      -- 
    ack_2704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nLSTATE_1380_1368_buf_ack_0, ack => nicRxFromMacDaemon_CP_2536_elements(33)); -- 
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_nLSTATE_1368_update_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_nLSTATE_1368_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_nLSTATE_1368_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_nLSTATE_1368_Update/ack
      -- 
    ack_2709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nLSTATE_1380_1368_buf_ack_1, ack => nicRxFromMacDaemon_CP_2536_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_S0_1369_sample_start__ps
      -- CP-element group 35: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_S0_1369_sample_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_S0_1369_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_S0_1369_sample_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_2536_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (2) 
      -- CP-element group 36: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_S0_1369_update_start__ps
      -- CP-element group 36: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_S0_1369_update_start_
      -- 
    -- Element group nicRxFromMacDaemon_CP_2536_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	38 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_S0_1369_update_completed__ps
      -- 
    nicRxFromMacDaemon_CP_2536_elements(37) <= nicRxFromMacDaemon_CP_2536_elements(38);
    -- CP-element group 38:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	37 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/R_S0_1369_update_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_2536_elements(38) is a control-delay.
    cp_element_38_delay: control_delay_element  generic map(name => " 38_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_2536_elements(36), ack => nicRxFromMacDaemon_CP_2536_elements(38), clk => clk, reset =>reset);
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	16 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	46 
    -- CP-element group 39: 	52 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	20 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1370_update_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2536_elements(16) & nicRxFromMacDaemon_CP_2536_elements(46) & nicRxFromMacDaemon_CP_2536_elements(52);
      gj_nicRxFromMacDaemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2536_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	18 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	43 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/RPIPE_mac_to_nic_data_1372_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/RPIPE_mac_to_nic_data_1372_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/RPIPE_mac_to_nic_data_1372_Sample/rr
      -- 
    rr_2730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2536_elements(40), ack => RPIPE_mac_to_nic_data_1372_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2536_elements(18) & nicRxFromMacDaemon_CP_2536_elements(43);
      gj_nicRxFromMacDaemon_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2536_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	42 
    -- CP-element group 41: 	20 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/RPIPE_mac_to_nic_data_1372_update_start_
      -- CP-element group 41: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/RPIPE_mac_to_nic_data_1372_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/RPIPE_mac_to_nic_data_1372_Update/cr
      -- 
    cr_2735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2536_elements(41), ack => RPIPE_mac_to_nic_data_1372_inst_req_1); -- 
    nicRxFromMacDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2536_elements(42) & nicRxFromMacDaemon_CP_2536_elements(20);
      gj_nicRxFromMacDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2536_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: 	19 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/RPIPE_mac_to_nic_data_1372_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/RPIPE_mac_to_nic_data_1372_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/RPIPE_mac_to_nic_data_1372_Sample/ra
      -- 
    ra_2731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mac_to_nic_data_1372_inst_ack_0, ack => nicRxFromMacDaemon_CP_2536_elements(42)); -- 
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43: 	21 
    -- CP-element group 43: 	51 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	40 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/phi_stmt_1370_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/RPIPE_mac_to_nic_data_1372_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/RPIPE_mac_to_nic_data_1372_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/RPIPE_mac_to_nic_data_1372_Update/ca
      -- 
    ca_2736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mac_to_nic_data_1372_inst_ack_1, ack => nicRxFromMacDaemon_CP_2536_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: 	25 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/MUX_1400_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/MUX_1400_start/$entry
      -- CP-element group 44: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/MUX_1400_start/req
      -- 
    req_2744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2536_elements(44), ack => MUX_1400_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2536_elements(43) & nicRxFromMacDaemon_CP_2536_elements(25) & nicRxFromMacDaemon_CP_2536_elements(46);
      gj_nicRxFromMacDaemon_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2536_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	47 
    -- CP-element group 45: 	49 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/MUX_1400_update_start_
      -- CP-element group 45: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/MUX_1400_complete/$entry
      -- CP-element group 45: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/MUX_1400_complete/req
      -- 
    req_2749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2536_elements(45), ack => MUX_1400_inst_req_1); -- 
    nicRxFromMacDaemon_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2536_elements(47) & nicRxFromMacDaemon_CP_2536_elements(49);
      gj_nicRxFromMacDaemon_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2536_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	39 
    -- CP-element group 46: 	44 
    -- CP-element group 46: 	23 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/MUX_1400_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/MUX_1400_start/$exit
      -- CP-element group 46: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/MUX_1400_start/ack
      -- 
    ack_2745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1400_inst_ack_0, ack => nicRxFromMacDaemon_CP_2536_elements(46)); -- 
    -- CP-element group 47:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: marked-successors 
    -- CP-element group 47: 	45 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/MUX_1400_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/MUX_1400_complete/$exit
      -- CP-element group 47: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/MUX_1400_complete/ack
      -- 
    ack_2750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1400_inst_ack_1, ack => nicRxFromMacDaemon_CP_2536_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	25 
    -- CP-element group 48: 	47 
    -- CP-element group 48: marked-predecessors 
    -- CP-element group 48: 	50 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_header_1391_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_header_1391_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_header_1391_Sample/req
      -- 
    req_2758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2536_elements(48), ack => WPIPE_nic_rx_to_header_1391_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2536_elements(25) & nicRxFromMacDaemon_CP_2536_elements(47) & nicRxFromMacDaemon_CP_2536_elements(50);
      gj_nicRxFromMacDaemon_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2536_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	45 
    -- CP-element group 49: 	23 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_header_1391_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_header_1391_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_header_1391_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_header_1391_Sample/ack
      -- CP-element group 49: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_header_1391_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_header_1391_Update/req
      -- 
    ack_2759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_header_1391_inst_ack_0, ack => nicRxFromMacDaemon_CP_2536_elements(49)); -- 
    req_2763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2536_elements(49), ack => WPIPE_nic_rx_to_header_1391_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	55 
    -- CP-element group 50: marked-successors 
    -- CP-element group 50: 	48 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_header_1391_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_header_1391_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_header_1391_Update/ack
      -- 
    ack_2764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_header_1391_inst_ack_1, ack => nicRxFromMacDaemon_CP_2536_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	43 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	53 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_packet_1402_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_packet_1402_Sample/req
      -- CP-element group 51: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_packet_1402_sample_start_
      -- 
    req_2772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2536_elements(51), ack => WPIPE_nic_rx_to_packet_1402_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2536_elements(43) & nicRxFromMacDaemon_CP_2536_elements(53);
      gj_nicRxFromMacDaemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2536_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	39 
    -- CP-element group 52:  members (6) 
      -- CP-element group 52: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_packet_1402_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_packet_1402_Sample/ack
      -- CP-element group 52: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_packet_1402_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_packet_1402_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_packet_1402_Update/req
      -- CP-element group 52: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_packet_1402_update_start_
      -- 
    ack_2773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_packet_1402_inst_ack_0, ack => nicRxFromMacDaemon_CP_2536_elements(52)); -- 
    req_2777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2536_elements(52), ack => WPIPE_nic_rx_to_packet_1402_inst_req_1); -- 
    -- CP-element group 53:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: marked-successors 
    -- CP-element group 53: 	51 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_packet_1402_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_packet_1402_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/WPIPE_nic_rx_to_packet_1402_Update/ack
      -- 
    ack_2778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_packet_1402_inst_ack_1, ack => nicRxFromMacDaemon_CP_2536_elements(53)); -- 
    -- CP-element group 54:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	16 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	17 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group nicRxFromMacDaemon_CP_2536_elements(54) is a control-delay.
    cp_element_54_delay: control_delay_element  generic map(name => " 54_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_2536_elements(16), ack => nicRxFromMacDaemon_CP_2536_elements(54), clk => clk, reset =>reset);
    -- CP-element group 55:  join  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	19 
    -- CP-element group 55: 	50 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	13 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_1333/do_while_stmt_1364/do_while_stmt_1364_loop_body/$exit
      -- 
    nicRxFromMacDaemon_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2536_elements(19) & nicRxFromMacDaemon_CP_2536_elements(50) & nicRxFromMacDaemon_CP_2536_elements(53);
      gj_nicRxFromMacDaemon_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2536_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	12 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_1333/do_while_stmt_1364/loop_exit/$exit
      -- CP-element group 56: 	 branch_block_stmt_1333/do_while_stmt_1364/loop_exit/ack
      -- 
    ack_2783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1364_branch_ack_0, ack => nicRxFromMacDaemon_CP_2536_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	12 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_1333/do_while_stmt_1364/loop_taken/$exit
      -- CP-element group 57: 	 branch_block_stmt_1333/do_while_stmt_1364/loop_taken/ack
      -- 
    ack_2787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1364_branch_ack_1, ack => nicRxFromMacDaemon_CP_2536_elements(57)); -- 
    -- CP-element group 58:  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	10 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	2 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1333/do_while_stmt_1364/$exit
      -- 
    nicRxFromMacDaemon_CP_2536_elements(58) <= nicRxFromMacDaemon_CP_2536_elements(10);
    -- CP-element group 59:  merge  fork  transition  place  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: 	2 
    -- CP-element group 59: 	5 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	3 
    -- CP-element group 59: 	4 
    -- CP-element group 59:  members (13) 
      -- CP-element group 59: 	 branch_block_stmt_1333/merge_stmt_1335_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_1333/merge_stmt_1335_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_1333/merge_stmt_1335_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_1333/merge_stmt_1335_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_1333/merge_stmt_1335__exit__
      -- CP-element group 59: 	 branch_block_stmt_1333/call_stmt_1345__entry__
      -- CP-element group 59: 	 branch_block_stmt_1333/call_stmt_1345/$entry
      -- CP-element group 59: 	 branch_block_stmt_1333/call_stmt_1345/call_stmt_1345_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_1333/call_stmt_1345/call_stmt_1345_update_start_
      -- CP-element group 59: 	 branch_block_stmt_1333/call_stmt_1345/call_stmt_1345_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1333/call_stmt_1345/call_stmt_1345_Sample/crr
      -- CP-element group 59: 	 branch_block_stmt_1333/call_stmt_1345/call_stmt_1345_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1333/call_stmt_1345/call_stmt_1345_Update/ccr
      -- 
    crr_2565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2536_elements(59), ack => call_stmt_1345_call_req_0); -- 
    ccr_2570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2536_elements(59), ack => call_stmt_1345_call_req_1); -- 
    nicRxFromMacDaemon_CP_2536_elements(59) <= OrReduce(nicRxFromMacDaemon_CP_2536_elements(0) & nicRxFromMacDaemon_CP_2536_elements(2) & nicRxFromMacDaemon_CP_2536_elements(5));
    nicRxFromMacDaemon_do_while_stmt_1364_terminator_2788: loop_terminator -- 
      generic map (name => " nicRxFromMacDaemon_do_while_stmt_1364_terminator_2788", max_iterations_in_flight =>7) 
      port map(loop_body_exit => nicRxFromMacDaemon_CP_2536_elements(13),loop_continue => nicRxFromMacDaemon_CP_2536_elements(57),loop_terminate => nicRxFromMacDaemon_CP_2536_elements(56),loop_back => nicRxFromMacDaemon_CP_2536_elements(11),loop_exit => nicRxFromMacDaemon_CP_2536_elements(10),clk => clk, reset => reset); -- 
    phi_stmt_1366_phi_seq_2718_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= nicRxFromMacDaemon_CP_2536_elements(26);
      nicRxFromMacDaemon_CP_2536_elements(31)<= src_sample_reqs(0);
      src_sample_acks(0)  <= nicRxFromMacDaemon_CP_2536_elements(33);
      nicRxFromMacDaemon_CP_2536_elements(32)<= src_update_reqs(0);
      src_update_acks(0)  <= nicRxFromMacDaemon_CP_2536_elements(34);
      nicRxFromMacDaemon_CP_2536_elements(27) <= phi_mux_reqs(0);
      triggers(1)  <= nicRxFromMacDaemon_CP_2536_elements(28);
      nicRxFromMacDaemon_CP_2536_elements(35)<= src_sample_reqs(1);
      src_sample_acks(1)  <= nicRxFromMacDaemon_CP_2536_elements(35);
      nicRxFromMacDaemon_CP_2536_elements(36)<= src_update_reqs(1);
      src_update_acks(1)  <= nicRxFromMacDaemon_CP_2536_elements(37);
      nicRxFromMacDaemon_CP_2536_elements(29) <= phi_mux_reqs(1);
      phi_stmt_1366_phi_seq_2718 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1366_phi_seq_2718") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => nicRxFromMacDaemon_CP_2536_elements(18), 
          phi_sample_ack => nicRxFromMacDaemon_CP_2536_elements(24), 
          phi_update_req => nicRxFromMacDaemon_CP_2536_elements(20), 
          phi_update_ack => nicRxFromMacDaemon_CP_2536_elements(25), 
          phi_mux_ack => nicRxFromMacDaemon_CP_2536_elements(30), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2670_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= nicRxFromMacDaemon_CP_2536_elements(14);
        preds(1)  <= nicRxFromMacDaemon_CP_2536_elements(15);
        entry_tmerge_2670 : transition_merge -- 
          generic map(name => " entry_tmerge_2670")
          port map (preds => preds, symbol_out => nicRxFromMacDaemon_CP_2536_elements(16));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_1349_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_1411_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u65_u73_1398_wire : std_logic_vector(72 downto 0);
    signal EQ_u2_u1_1384_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1387_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1394_wire : std_logic_vector(0 downto 0);
    signal LSTATE_1366 : std_logic_vector(1 downto 0);
    signal MUX_1400_wire : std_logic_vector(72 downto 0);
    signal NOT_u1_u1_1350_wire : std_logic_vector(0 downto 0);
    signal NOT_u4_u4_1340_wire_constant : std_logic_vector(3 downto 0);
    signal NOT_u4_u4_1358_wire_constant : std_logic_vector(3 downto 0);
    signal RPIPE_CONTROL_REGISTER_1347_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CONTROL_REGISTER_1409_wire : std_logic_vector(31 downto 0);
    signal RPIPE_mac_to_nic_data_1372_wire : std_logic_vector(72 downto 0);
    signal RX_1370 : std_logic_vector(72 downto 0);
    signal R_HEADER_TKEEP_1397_wire_constant : std_logic_vector(7 downto 0);
    signal R_S0_1369_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_1383_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_1386_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_1393_wire_constant : std_logic_vector(1 downto 0);
    signal ignore_resp0_1345 : std_logic_vector(31 downto 0);
    signal ignore_resp1_1363 : std_logic_vector(31 downto 0);
    signal konst_1341_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1348_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1359_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1410_wire_constant : std_logic_vector(31 downto 0);
    signal nLSTATE_1380 : std_logic_vector(1 downto 0);
    signal nLSTATE_1380_1368_buffered : std_logic_vector(1 downto 0);
    signal slice_1396_wire : std_logic_vector(64 downto 0);
    signal type_cast_1337_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1343_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1355_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1361_wire_constant : std_logic_vector(31 downto 0);
    signal write_to_header_1389 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_1340_wire_constant <= "1111";
    NOT_u4_u4_1358_wire_constant <= "1111";
    R_HEADER_TKEEP_1397_wire_constant <= "00111111";
    R_S0_1369_wire_constant <= "00";
    R_S0_1383_wire_constant <= "00";
    R_S1_1386_wire_constant <= "01";
    R_S1_1393_wire_constant <= "01";
    konst_1341_wire_constant <= "010110";
    konst_1348_wire_constant <= "00000000000000000000000000000000";
    konst_1359_wire_constant <= "010110";
    konst_1410_wire_constant <= "00000000000000000000000000000000";
    type_cast_1337_wire_constant <= "0";
    type_cast_1343_wire_constant <= "00000000000000000000000000000000";
    type_cast_1355_wire_constant <= "0";
    type_cast_1361_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_1366: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nLSTATE_1380_1368_buffered & R_S0_1369_wire_constant;
      req <= phi_stmt_1366_req_0 & phi_stmt_1366_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1366",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1366_ack_0,
          idata => idata,
          odata => LSTATE_1366,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1366
    MUX_1400_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      signal sample_req_ug, sample_ack_ug, update_req_ug, update_ack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      sample_req_ug(0) <= MUX_1400_inst_req_0;
      MUX_1400_inst_ack_0<= sample_ack_ug(0);
      update_req_ug(0) <= MUX_1400_inst_req_1;
      MUX_1400_inst_ack_1<= update_ack_ug(0);
      guard_vector(0) <=  write_to_header_1389(0);
      MUX_1400_inst_gI: SplitGuardInterface generic map(name => "MUX_1400_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_ug,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_ug,
        cr_in => update_req_ug,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_ug,
        guards => guard_vector); -- 
      MUX_1400_inst: SelectSplitProtocol generic map(name => "MUX_1400_inst", data_width => 73, buffering => 1, flow_through => false, full_rate => true) -- 
        port map( x => CONCAT_u65_u73_1398_wire, y => RX_1370, sel => EQ_u2_u1_1394_wire, z => MUX_1400_wire, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through slice operator slice_1396_inst
    slice_1396_wire <= RX_1370(72 downto 8);
    nLSTATE_1380_1368_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nLSTATE_1380_1368_buf_req_0;
      nLSTATE_1380_1368_buf_ack_0<= wack(0);
      rreq(0) <= nLSTATE_1380_1368_buf_req_1;
      nLSTATE_1380_1368_buf_ack_1<= rack(0);
      nLSTATE_1380_1368_buf : InterlockBuffer generic map ( -- 
        name => "nLSTATE_1380_1368_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nLSTATE_1380,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nLSTATE_1380_1368_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1370
    process(RPIPE_mac_to_nic_data_1372_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_mac_to_nic_data_1372_wire(72 downto 0);
      RX_1370 <= tmp_var; -- 
    end process;
    do_while_stmt_1364_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_1411_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1364_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1364_branch_req_0,
          ack0 => do_while_stmt_1364_branch_ack_0,
          ack1 => do_while_stmt_1364_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1346_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1350_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1346_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1346_branch_req_0,
          ack0 => if_stmt_1346_branch_ack_0,
          ack1 => if_stmt_1346_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator BITSEL_u32_u1_1349_inst
    process(RPIPE_CONTROL_REGISTER_1347_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1347_wire, konst_1348_wire_constant, tmp_var);
      BITSEL_u32_u1_1349_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1411_inst
    process(RPIPE_CONTROL_REGISTER_1409_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1409_wire, konst_1410_wire_constant, tmp_var);
      BITSEL_u32_u1_1411_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u65_u73_1398_inst
    process(slice_1396_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1396_wire, R_HEADER_TKEEP_1397_wire_constant, tmp_var);
      CONCAT_u65_u73_1398_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1384_inst
    process(LSTATE_1366) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_1366, R_S0_1383_wire_constant, tmp_var);
      EQ_u2_u1_1384_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1387_inst
    process(LSTATE_1366) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_1366, R_S1_1386_wire_constant, tmp_var);
      EQ_u2_u1_1387_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1394_inst
    process(LSTATE_1366) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_1366, R_S1_1393_wire_constant, tmp_var);
      EQ_u2_u1_1394_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1350_inst
    process(BITSEL_u32_u1_1349_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_1349_wire, tmp_var);
      NOT_u1_u1_1350_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1388_inst
    process(EQ_u2_u1_1384_wire, EQ_u2_u1_1387_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u2_u1_1384_wire, EQ_u2_u1_1387_wire, tmp_var);
      write_to_header_1389 <= tmp_var; --
    end process;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1347_wire <= CONTROL_REGISTER;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1409_wire <= CONTROL_REGISTER;
    -- shared inport operator group (2) : RPIPE_mac_to_nic_data_1372_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_mac_to_nic_data_1372_inst_req_0;
      RPIPE_mac_to_nic_data_1372_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_mac_to_nic_data_1372_inst_req_1;
      RPIPE_mac_to_nic_data_1372_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_mac_to_nic_data_1372_wire <= data_out(72 downto 0);
      mac_to_nic_data_read_2_gI: SplitGuardInterface generic map(name => "mac_to_nic_data_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      mac_to_nic_data_read_2: InputPortRevised -- 
        generic map ( name => "mac_to_nic_data_read_2", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => mac_to_nic_data_pipe_read_req(0),
          oack => mac_to_nic_data_pipe_read_ack(0),
          odata => mac_to_nic_data_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared outport operator group (0) : WPIPE_nic_rx_to_header_1391_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_rx_to_header_1391_inst_req_0;
      WPIPE_nic_rx_to_header_1391_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_rx_to_header_1391_inst_req_1;
      WPIPE_nic_rx_to_header_1391_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_to_header_1389(0);
      data_in <= MUX_1400_wire;
      nic_rx_to_header_write_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_header_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_header_write_0: OutputPortRevised -- 
        generic map ( name => "nic_rx_to_header", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_rx_to_header_pipe_write_req(0),
          oack => nic_rx_to_header_pipe_write_ack(0),
          odata => nic_rx_to_header_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_nic_rx_to_packet_1402_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_rx_to_packet_1402_inst_req_0;
      WPIPE_nic_rx_to_packet_1402_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_rx_to_packet_1402_inst_req_1;
      WPIPE_nic_rx_to_packet_1402_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= RX_1370;
      nic_rx_to_packet_write_1_gI: SplitGuardInterface generic map(name => "nic_rx_to_packet_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_packet_write_1: OutputPortRevised -- 
        generic map ( name => "nic_rx_to_packet", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_rx_to_packet_pipe_write_req(0),
          oack => nic_rx_to_packet_pipe_write_ack(0),
          odata => nic_rx_to_packet_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_1363_call call_stmt_1345_call 
    AccessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(85 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1363_call_req_0;
      reqL_unguarded(0) <= call_stmt_1345_call_req_0;
      call_stmt_1363_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1345_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1363_call_req_1;
      reqR_unguarded(0) <= call_stmt_1345_call_req_1;
      call_stmt_1363_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1345_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      AccessRegister_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "AccessRegister_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      AccessRegister_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "AccessRegister_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      AccessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1355_wire_constant & NOT_u4_u4_1358_wire_constant & konst_1359_wire_constant & type_cast_1361_wire_constant & type_cast_1337_wire_constant & NOT_u4_u4_1340_wire_constant & konst_1341_wire_constant & type_cast_1343_wire_constant;
      ignore_resp1_1363 <= data_out(63 downto 32);
      ignore_resp0_1345 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 86,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    volatile_operator_nextLSTATE_3876: nextLSTATE_Volatile port map(RX => RX_1370, LSTATE => LSTATE_1366, nLSTATE => nLSTATE_1380); 
    -- 
  end Block; -- data_path
  -- 
end nicRxFromMacDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity popFromQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    lock : in  std_logic_vector(0 downto 0);
    q_base_address : in  std_logic_vector(35 downto 0);
    q_r_data : out  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
    setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
    releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
    releaseMutex_call_data : out  std_logic_vector(35 downto 0);
    releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
    releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
    releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
    releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
    getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
    getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
    getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
    getQueueElement_call_data : out  std_logic_vector(67 downto 0);
    getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
    getQueueElement_return_data : in   std_logic_vector(31 downto 0);
    getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
    acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
    acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
    acquireMutex_call_data : out  std_logic_vector(35 downto 0);
    acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
    acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
    acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
    acquireMutex_return_data : in   std_logic_vector(0 downto 0);
    acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity popFromQueue;
architecture popFromQueue_arch of popFromQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 37)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 33)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal q_r_data_buffer :  std_logic_vector(31 downto 0);
  signal q_r_data_update_enable: Boolean;
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal popFromQueue_CP_604_start: Boolean;
  signal popFromQueue_CP_604_symbol: Boolean;
  -- volatile/operator module components. 
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component releaseMutex is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      read_pointer : in  std_logic_vector(31 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component acquireMutex is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_492_call_req_0 : boolean;
  signal call_stmt_522_call_req_0 : boolean;
  signal call_stmt_522_call_ack_0 : boolean;
  signal call_stmt_522_call_req_1 : boolean;
  signal call_stmt_522_call_ack_1 : boolean;
  signal call_stmt_497_call_req_0 : boolean;
  signal call_stmt_497_call_ack_0 : boolean;
  signal call_stmt_492_call_ack_0 : boolean;
  signal call_stmt_492_call_req_1 : boolean;
  signal call_stmt_527_call_req_0 : boolean;
  signal call_stmt_527_call_ack_0 : boolean;
  signal call_stmt_527_call_req_1 : boolean;
  signal call_stmt_527_call_ack_1 : boolean;
  signal call_stmt_492_call_ack_1 : boolean;
  signal call_stmt_497_call_req_1 : boolean;
  signal call_stmt_497_call_ack_1 : boolean;
  signal call_stmt_538_call_req_0 : boolean;
  signal call_stmt_538_call_ack_0 : boolean;
  signal call_stmt_538_call_req_1 : boolean;
  signal call_stmt_538_call_ack_1 : boolean;
  signal W_status_539_inst_req_0 : boolean;
  signal W_status_539_inst_ack_0 : boolean;
  signal W_status_539_inst_req_1 : boolean;
  signal W_status_539_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "popFromQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 37) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= lock;
  lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(36 downto 1) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(36 downto 1);
  in_buffer_data_in(tag_length + 36 downto 37) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 36 downto 37);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  popFromQueue_CP_604_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "popFromQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 33) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= q_r_data_buffer;
  q_r_data <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(32 downto 32) <= status_buffer;
  status <= out_buffer_data_out(32 downto 32);
  out_buffer_data_in(tag_length + 32 downto 33) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 32 downto 33);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= popFromQueue_CP_604_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= popFromQueue_CP_604_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= popFromQueue_CP_604_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  popFromQueue_CP_604: Block -- control-path 
    signal popFromQueue_CP_604_elements: BooleanArray(14 downto 0);
    -- 
  begin -- 
    popFromQueue_CP_604_elements(0) <= popFromQueue_CP_604_start;
    popFromQueue_CP_604_symbol <= popFromQueue_CP_604_elements(14);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_492/call_stmt_492_sample_start_
      -- CP-element group 0: 	 call_stmt_492/call_stmt_492_Sample/$entry
      -- CP-element group 0: 	 call_stmt_492/call_stmt_492_Sample/crr
      -- CP-element group 0: 	 call_stmt_492/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_492/call_stmt_492_Update/$entry
      -- CP-element group 0: 	 call_stmt_492/call_stmt_492_Update/ccr
      -- CP-element group 0: 	 call_stmt_492/call_stmt_492_update_start_
      -- 
    crr_617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_604_elements(0), ack => call_stmt_492_call_req_0); -- 
    ccr_622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_604_elements(0), ack => call_stmt_492_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_492/call_stmt_492_Sample/$exit
      -- CP-element group 1: 	 call_stmt_492/call_stmt_492_Sample/cra
      -- CP-element group 1: 	 call_stmt_492/call_stmt_492_sample_completed_
      -- 
    cra_618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_492_call_ack_0, ack => popFromQueue_CP_604_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	9 
    -- CP-element group 2:  members (17) 
      -- CP-element group 2: 	 call_stmt_492/$exit
      -- CP-element group 2: 	 call_stmt_492/call_stmt_492_update_completed_
      -- CP-element group 2: 	 call_stmt_497_to_call_stmt_527/call_stmt_522_Update/$entry
      -- CP-element group 2: 	 call_stmt_497_to_call_stmt_527/call_stmt_522_Update/ccr
      -- CP-element group 2: 	 call_stmt_497_to_call_stmt_527/call_stmt_497_Sample/$entry
      -- CP-element group 2: 	 call_stmt_497_to_call_stmt_527/call_stmt_497_Sample/crr
      -- CP-element group 2: 	 call_stmt_497_to_call_stmt_527/call_stmt_497_Update/$entry
      -- CP-element group 2: 	 call_stmt_492/call_stmt_492_Update/$exit
      -- CP-element group 2: 	 call_stmt_497_to_call_stmt_527/call_stmt_527_update_start_
      -- CP-element group 2: 	 call_stmt_497_to_call_stmt_527/call_stmt_527_Update/$entry
      -- CP-element group 2: 	 call_stmt_497_to_call_stmt_527/call_stmt_527_Update/ccr
      -- CP-element group 2: 	 call_stmt_497_to_call_stmt_527/call_stmt_497_update_start_
      -- CP-element group 2: 	 call_stmt_497_to_call_stmt_527/$entry
      -- CP-element group 2: 	 call_stmt_497_to_call_stmt_527/call_stmt_497_sample_start_
      -- CP-element group 2: 	 call_stmt_492/call_stmt_492_Update/cca
      -- CP-element group 2: 	 call_stmt_497_to_call_stmt_527/call_stmt_497_Update/ccr
      -- CP-element group 2: 	 call_stmt_497_to_call_stmt_527/call_stmt_522_update_start_
      -- 
    cca_623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_492_call_ack_1, ack => popFromQueue_CP_604_elements(2)); -- 
    crr_634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_604_elements(2), ack => call_stmt_497_call_req_0); -- 
    ccr_639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_604_elements(2), ack => call_stmt_497_call_req_1); -- 
    ccr_653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_604_elements(2), ack => call_stmt_522_call_req_1); -- 
    ccr_667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_604_elements(2), ack => call_stmt_527_call_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_497_to_call_stmt_527/call_stmt_497_Sample/$exit
      -- CP-element group 3: 	 call_stmt_497_to_call_stmt_527/call_stmt_497_Sample/cra
      -- CP-element group 3: 	 call_stmt_497_to_call_stmt_527/call_stmt_497_sample_completed_
      -- 
    cra_635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_497_call_ack_0, ack => popFromQueue_CP_604_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 call_stmt_497_to_call_stmt_527/call_stmt_522_Sample/$entry
      -- CP-element group 4: 	 call_stmt_497_to_call_stmt_527/call_stmt_522_Sample/crr
      -- CP-element group 4: 	 call_stmt_497_to_call_stmt_527/call_stmt_497_Update/$exit
      -- CP-element group 4: 	 call_stmt_497_to_call_stmt_527/call_stmt_497_update_completed_
      -- CP-element group 4: 	 call_stmt_497_to_call_stmt_527/call_stmt_497_Update/cca
      -- CP-element group 4: 	 call_stmt_497_to_call_stmt_527/call_stmt_522_sample_start_
      -- 
    cca_640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_497_call_ack_1, ack => popFromQueue_CP_604_elements(4)); -- 
    crr_648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_604_elements(4), ack => call_stmt_522_call_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_497_to_call_stmt_527/call_stmt_522_Sample/$exit
      -- CP-element group 5: 	 call_stmt_497_to_call_stmt_527/call_stmt_522_Sample/cra
      -- CP-element group 5: 	 call_stmt_497_to_call_stmt_527/call_stmt_522_sample_completed_
      -- 
    cra_649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_522_call_ack_0, ack => popFromQueue_CP_604_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 call_stmt_497_to_call_stmt_527/call_stmt_522_Update/$exit
      -- CP-element group 6: 	 call_stmt_497_to_call_stmt_527/call_stmt_522_Update/cca
      -- CP-element group 6: 	 call_stmt_497_to_call_stmt_527/call_stmt_522_update_completed_
      -- 
    cca_654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_522_call_ack_1, ack => popFromQueue_CP_604_elements(6)); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_497_to_call_stmt_527/call_stmt_527_sample_start_
      -- CP-element group 7: 	 call_stmt_497_to_call_stmt_527/call_stmt_527_Sample/$entry
      -- CP-element group 7: 	 call_stmt_497_to_call_stmt_527/call_stmt_527_Sample/crr
      -- 
    crr_662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_604_elements(7), ack => call_stmt_527_call_req_0); -- 
    popFromQueue_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "popFromQueue_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= popFromQueue_CP_604_elements(4) & popFromQueue_CP_604_elements(6);
      gj_popFromQueue_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_604_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_497_to_call_stmt_527/call_stmt_527_sample_completed_
      -- CP-element group 8: 	 call_stmt_497_to_call_stmt_527/call_stmt_527_Sample/$exit
      -- CP-element group 8: 	 call_stmt_497_to_call_stmt_527/call_stmt_527_Sample/cra
      -- 
    cra_663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_527_call_ack_0, ack => popFromQueue_CP_604_elements(8)); -- 
    -- CP-element group 9:  fork  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9:  members (17) 
      -- CP-element group 9: 	 call_stmt_497_to_call_stmt_527/call_stmt_527_update_completed_
      -- CP-element group 9: 	 call_stmt_497_to_call_stmt_527/call_stmt_527_Update/$exit
      -- CP-element group 9: 	 call_stmt_497_to_call_stmt_527/call_stmt_527_Update/cca
      -- CP-element group 9: 	 call_stmt_538_to_assign_stmt_541/$entry
      -- CP-element group 9: 	 call_stmt_538_to_assign_stmt_541/call_stmt_538_sample_start_
      -- CP-element group 9: 	 call_stmt_497_to_call_stmt_527/$exit
      -- CP-element group 9: 	 call_stmt_538_to_assign_stmt_541/call_stmt_538_update_start_
      -- CP-element group 9: 	 call_stmt_538_to_assign_stmt_541/call_stmt_538_Sample/$entry
      -- CP-element group 9: 	 call_stmt_538_to_assign_stmt_541/call_stmt_538_Sample/crr
      -- CP-element group 9: 	 call_stmt_538_to_assign_stmt_541/call_stmt_538_Update/$entry
      -- CP-element group 9: 	 call_stmt_538_to_assign_stmt_541/call_stmt_538_Update/ccr
      -- CP-element group 9: 	 call_stmt_538_to_assign_stmt_541/assign_stmt_541_sample_start_
      -- CP-element group 9: 	 call_stmt_538_to_assign_stmt_541/assign_stmt_541_update_start_
      -- CP-element group 9: 	 call_stmt_538_to_assign_stmt_541/assign_stmt_541_Sample/$entry
      -- CP-element group 9: 	 call_stmt_538_to_assign_stmt_541/assign_stmt_541_Sample/req
      -- CP-element group 9: 	 call_stmt_538_to_assign_stmt_541/assign_stmt_541_Update/$entry
      -- CP-element group 9: 	 call_stmt_538_to_assign_stmt_541/assign_stmt_541_Update/req
      -- 
    cca_668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_527_call_ack_1, ack => popFromQueue_CP_604_elements(9)); -- 
    crr_679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_604_elements(9), ack => call_stmt_538_call_req_0); -- 
    ccr_684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_604_elements(9), ack => call_stmt_538_call_req_1); -- 
    req_693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_604_elements(9), ack => W_status_539_inst_req_0); -- 
    req_698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_604_elements(9), ack => W_status_539_inst_req_1); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_538_to_assign_stmt_541/call_stmt_538_sample_completed_
      -- CP-element group 10: 	 call_stmt_538_to_assign_stmt_541/call_stmt_538_Sample/$exit
      -- CP-element group 10: 	 call_stmt_538_to_assign_stmt_541/call_stmt_538_Sample/cra
      -- 
    cra_680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_538_call_ack_0, ack => popFromQueue_CP_604_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_538_to_assign_stmt_541/call_stmt_538_update_completed_
      -- CP-element group 11: 	 call_stmt_538_to_assign_stmt_541/call_stmt_538_Update/$exit
      -- CP-element group 11: 	 call_stmt_538_to_assign_stmt_541/call_stmt_538_Update/cca
      -- 
    cca_685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_538_call_ack_1, ack => popFromQueue_CP_604_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_538_to_assign_stmt_541/assign_stmt_541_sample_completed_
      -- CP-element group 12: 	 call_stmt_538_to_assign_stmt_541/assign_stmt_541_Sample/$exit
      -- CP-element group 12: 	 call_stmt_538_to_assign_stmt_541/assign_stmt_541_Sample/ack
      -- 
    ack_694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_status_539_inst_ack_0, ack => popFromQueue_CP_604_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_538_to_assign_stmt_541/assign_stmt_541_update_completed_
      -- CP-element group 13: 	 call_stmt_538_to_assign_stmt_541/assign_stmt_541_Update/$exit
      -- CP-element group 13: 	 call_stmt_538_to_assign_stmt_541/assign_stmt_541_Update/ack
      -- 
    ack_699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_status_539_inst_ack_1, ack => popFromQueue_CP_604_elements(13)); -- 
    -- CP-element group 14:  join  transition  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 $exit
      -- CP-element group 14: 	 call_stmt_538_to_assign_stmt_541/$exit
      -- 
    popFromQueue_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "popFromQueue_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= popFromQueue_CP_604_elements(11) & popFromQueue_CP_604_elements(13);
      gj_popFromQueue_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_604_elements(14), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_515_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_507_wire_constant : std_logic_vector(31 downto 0);
    signal konst_512_wire_constant : std_logic_vector(31 downto 0);
    signal konst_514_wire_constant : std_logic_vector(31 downto 0);
    signal m_ok_492 : std_logic_vector(0 downto 0);
    signal next_rp_517 : std_logic_vector(31 downto 0);
    signal q_empty_502 : std_logic_vector(0 downto 0);
    signal read_pointer_497 : std_logic_vector(31 downto 0);
    signal round_off_509 : std_logic_vector(0 downto 0);
    signal write_pointer_497 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    SUB_u32_u32_507_wire_constant <= "00000000000000000000000000000111";
    konst_512_wire_constant <= "00000000000000000000000000000000";
    konst_514_wire_constant <= "00000000000000000000000000000001";
    -- flow-through select operator MUX_516_inst
    next_rp_517 <= konst_512_wire_constant when (round_off_509(0) /=  '0') else ADD_u32_u32_515_wire;
    W_status_539_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_status_539_inst_req_0;
      W_status_539_inst_ack_0<= wack(0);
      rreq(0) <= W_status_539_inst_req_1;
      W_status_539_inst_ack_1<= rack(0);
      W_status_539_inst : InterlockBuffer generic map ( -- 
        name => "W_status_539_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => q_empty_502,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => status_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- binary operator ADD_u32_u32_515_inst
    process(read_pointer_497) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(read_pointer_497, konst_514_wire_constant, tmp_var);
      ADD_u32_u32_515_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_501_inst
    process(write_pointer_497, read_pointer_497) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(write_pointer_497, read_pointer_497, tmp_var);
      q_empty_502 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_508_inst
    process(read_pointer_497) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(read_pointer_497, SUB_u32_u32_507_wire_constant, tmp_var);
      round_off_509 <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_492_call 
    acquireMutex_call_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_492_call_req_0;
      call_stmt_492_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_492_call_req_1;
      call_stmt_492_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      acquireMutex_call_group_0_gI: SplitGuardInterface generic map(name => "acquireMutex_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      m_ok_492 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => acquireMutex_call_reqs(0),
          ackR => acquireMutex_call_acks(0),
          dataR => acquireMutex_call_data(35 downto 0),
          tagR => acquireMutex_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => acquireMutex_return_acks(0), -- cross-over
          ackL => acquireMutex_return_reqs(0), -- cross-over
          dataL => acquireMutex_return_data(0 downto 0),
          tagL => acquireMutex_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_497_call 
    getQueuePointers_call_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_497_call_req_0;
      call_stmt_497_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_497_call_req_1;
      call_stmt_497_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueuePointers_call_group_1_gI: SplitGuardInterface generic map(name => "getQueuePointers_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      write_pointer_497 <= data_out(63 downto 32);
      read_pointer_497 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueuePointers_call_reqs(0),
          ackR => getQueuePointers_call_acks(0),
          dataR => getQueuePointers_call_data(35 downto 0),
          tagR => getQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueuePointers_return_acks(0), -- cross-over
          ackL => getQueuePointers_return_reqs(0), -- cross-over
          dataL => getQueuePointers_return_data(63 downto 0),
          tagL => getQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_522_call 
    getQueueElement_call_group_2: Block -- 
      signal data_in: std_logic_vector(67 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_522_call_req_0;
      call_stmt_522_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_522_call_req_1;
      call_stmt_522_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_502(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueElement_call_group_2_gI: SplitGuardInterface generic map(name => "getQueueElement_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & read_pointer_497;
      q_r_data_buffer <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 68,
        owidth => 68,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueElement_call_reqs(0),
          ackR => getQueueElement_call_acks(0),
          dataR => getQueueElement_call_data(67 downto 0),
          tagR => getQueueElement_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueElement_return_acks(0), -- cross-over
          ackL => getQueueElement_return_reqs(0), -- cross-over
          dataL => getQueueElement_return_data(31 downto 0),
          tagL => getQueueElement_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_527_call 
    setQueuePointers_call_group_3: Block -- 
      signal data_in: std_logic_vector(99 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_527_call_req_0;
      call_stmt_527_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_527_call_req_1;
      call_stmt_527_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_502(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueuePointers_call_group_3_gI: SplitGuardInterface generic map(name => "setQueuePointers_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & write_pointer_497 & next_rp_517;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 100,
        owidth => 100,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueuePointers_call_reqs(0),
          ackR => setQueuePointers_call_acks(0),
          dataR => setQueuePointers_call_data(99 downto 0),
          tagR => setQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueuePointers_return_acks(0), -- cross-over
          ackL => setQueuePointers_return_reqs(0), -- cross-over
          tagL => setQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_538_call 
    releaseMutex_call_group_4: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_538_call_req_0;
      call_stmt_538_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_538_call_req_1;
      call_stmt_538_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      releaseMutex_call_group_4_gI: SplitGuardInterface generic map(name => "releaseMutex_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => releaseMutex_call_reqs(0),
          ackR => releaseMutex_call_acks(0),
          dataR => releaseMutex_call_data(35 downto 0),
          tagR => releaseMutex_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => releaseMutex_return_acks(0), -- cross-over
          ackL => releaseMutex_return_reqs(0), -- cross-over
          tagL => releaseMutex_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- 
  end Block; -- data_path
  -- 
end popFromQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity populateRxQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    rx_buffer_pointer : in  std_logic_vector(35 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
    NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity populateRxQueue;
architecture populateRxQueue_arch of populateRxQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rx_buffer_pointer_buffer :  std_logic_vector(35 downto 0);
  signal rx_buffer_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal populateRxQueue_CP_1330_start: Boolean;
  signal populateRxQueue_CP_1330_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component delay_time_Operator is -- 
    port ( -- 
      sample_req: in boolean;
      sample_ack: out boolean;
      update_req: in boolean;
      update_ack: out boolean;
      T : in  std_logic_vector(31 downto 0);
      delay_done : out  std_logic_vector(0 downto 0);
      clk, reset: in std_logic
      -- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_931_call_req_0 : boolean;
  signal call_stmt_931_call_req_1 : boolean;
  signal call_stmt_931_call_ack_0 : boolean;
  signal call_stmt_931_call_ack_1 : boolean;
  signal if_stmt_945_branch_ack_1 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_inst_ack_1 : boolean;
  signal if_stmt_945_branch_req_0 : boolean;
  signal if_stmt_951_branch_req_0 : boolean;
  signal call_stmt_914_call_req_0 : boolean;
  signal call_stmt_914_call_ack_0 : boolean;
  signal if_stmt_945_branch_ack_0 : boolean;
  signal if_stmt_951_branch_ack_0 : boolean;
  signal phi_stmt_883_req_1 : boolean;
  signal AND_u6_u6_892_inst_req_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_inst_req_1 : boolean;
  signal call_stmt_950_call_req_0 : boolean;
  signal call_stmt_914_call_ack_1 : boolean;
  signal AND_u6_u6_892_inst_ack_0 : boolean;
  signal AND_u6_u6_892_inst_ack_1 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_inst_req_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_inst_ack_0 : boolean;
  signal phi_stmt_883_req_0 : boolean;
  signal if_stmt_951_branch_ack_1 : boolean;
  signal call_stmt_914_call_req_1 : boolean;
  signal AND_u6_u6_892_inst_req_1 : boolean;
  signal AND_u6_u6_940_inst_ack_1 : boolean;
  signal AND_u6_u6_940_inst_req_1 : boolean;
  signal AND_u6_u6_940_inst_ack_0 : boolean;
  signal n_q_index_941_893_buf_ack_1 : boolean;
  signal call_stmt_950_call_ack_1 : boolean;
  signal call_stmt_950_call_req_1 : boolean;
  signal n_q_index_941_893_buf_req_1 : boolean;
  signal call_stmt_950_call_ack_0 : boolean;
  signal AND_u6_u6_940_inst_req_0 : boolean;
  signal phi_stmt_883_ack_0 : boolean;
  signal n_q_index_941_893_buf_ack_0 : boolean;
  signal n_q_index_941_893_buf_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "populateRxQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= rx_buffer_pointer;
  rx_buffer_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  populateRxQueue_CP_1330_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "populateRxQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= populateRxQueue_CP_1330_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= populateRxQueue_CP_1330_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= populateRxQueue_CP_1330_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  populateRxQueue_CP_1330: Block -- control-path 
    signal populateRxQueue_CP_1330_elements: BooleanArray(25 downto 0);
    -- 
  begin -- 
    populateRxQueue_CP_1330_elements(0) <= populateRxQueue_CP_1330_start;
    populateRxQueue_CP_1330_symbol <= populateRxQueue_CP_1330_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	17 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 branch_block_stmt_881/merge_stmt_882_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_881/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_881/merge_stmt_882__entry__
      -- CP-element group 0: 	 branch_block_stmt_881/branch_block_stmt_881__entry__
      -- 
    -- CP-element group 1:  merge  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	14 
    -- CP-element group 1: 	16 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_881/if_stmt_945__exit__
      -- CP-element group 1: 	 branch_block_stmt_881/$exit
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_881/branch_block_stmt_881__exit__
      -- 
    populateRxQueue_CP_1330_elements(1) <= OrReduce(populateRxQueue_CP_1330_elements(14) & populateRxQueue_CP_1330_elements(16));
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	25 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_914_Sample/cra
      -- CP-element group 2: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_914_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_914_sample_completed_
      -- 
    cra_1355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_914_call_ack_0, ack => populateRxQueue_CP_1330_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	25 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_931_Sample/crr
      -- CP-element group 3: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_931_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_914_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_931_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_914_Update/cca
      -- CP-element group 3: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_914_Update/$exit
      -- 
    cca_1360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_914_call_ack_1, ack => populateRxQueue_CP_1330_elements(3)); -- 
    crr_1368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1330_elements(3), ack => call_stmt_931_call_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_931_Sample/cra
      -- CP-element group 4: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_931_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_931_Sample/$exit
      -- 
    cra_1369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_931_call_ack_0, ack => populateRxQueue_CP_1330_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	25 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	8 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_931_Update/cca
      -- CP-element group 5: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_931_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_931_update_completed_
      -- 
    cca_1374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_931_call_ack_1, ack => populateRxQueue_CP_1330_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	25 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/AND_u6_u6_940_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/AND_u6_u6_940_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/AND_u6_u6_940_sample_completed_
      -- 
    ra_1383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_940_inst_ack_0, ack => populateRxQueue_CP_1330_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	25 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/AND_u6_u6_940_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/AND_u6_u6_940_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/AND_u6_u6_940_update_completed_
      -- 
    ca_1388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_940_inst_ack_1, ack => populateRxQueue_CP_1330_elements(7)); -- 
    -- CP-element group 8:  branch  join  transition  place  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	5 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (22) 
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945_else_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945_eval_test/NOT_u1_u1_947/SplitProtocol/Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945__entry__
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945_dead_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945_eval_test/branch_req
      -- CP-element group 8: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/$exit
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945_if_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945_eval_test/NOT_u1_u1_947/$entry
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945_eval_test/NOT_u1_u1_947/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945_eval_test/NOT_u1_u1_947/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941__exit__
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945_eval_test/$exit
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945_eval_test/$entry
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945_eval_test/NOT_u1_u1_947/SplitProtocol/$exit
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945_eval_test/NOT_u1_u1_947/$exit
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945_eval_test/NOT_u1_u1_947/SplitProtocol/Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945_eval_test/NOT_u1_u1_947/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945_eval_test/NOT_u1_u1_947/SplitProtocol/Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_881/NOT_u1_u1_947_place
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945_eval_test/NOT_u1_u1_947/SplitProtocol/Update/cr
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945_eval_test/NOT_u1_u1_947/SplitProtocol/Update/ca
      -- CP-element group 8: 	 branch_block_stmt_881/if_stmt_945_eval_test/NOT_u1_u1_947/SplitProtocol/Update/$entry
      -- 
    branch_req_1412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1330_elements(8), ack => if_stmt_945_branch_req_0); -- 
    populateRxQueue_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "populateRxQueue_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_1330_elements(5) & populateRxQueue_CP_1330_elements(7);
      gj_populateRxQueue_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_1330_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  fork  transition  place  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (10) 
      -- CP-element group 9: 	 branch_block_stmt_881/if_stmt_945_if_link/if_choice_transition
      -- CP-element group 9: 	 branch_block_stmt_881/call_stmt_950/call_stmt_950_update_start_
      -- CP-element group 9: 	 branch_block_stmt_881/call_stmt_950__entry__
      -- CP-element group 9: 	 branch_block_stmt_881/call_stmt_950/call_stmt_950_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_881/call_stmt_950/call_stmt_950_Sample/crr
      -- CP-element group 9: 	 branch_block_stmt_881/if_stmt_945_if_link/$exit
      -- CP-element group 9: 	 branch_block_stmt_881/call_stmt_950/$entry
      -- CP-element group 9: 	 branch_block_stmt_881/call_stmt_950/call_stmt_950_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_881/call_stmt_950/call_stmt_950_Update/ccr
      -- CP-element group 9: 	 branch_block_stmt_881/call_stmt_950/call_stmt_950_Update/$entry
      -- 
    if_choice_transition_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_945_branch_ack_1, ack => populateRxQueue_CP_1330_elements(9)); -- 
    crr_1436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1330_elements(9), ack => call_stmt_950_call_req_0); -- 
    ccr_1441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1330_elements(9), ack => call_stmt_950_call_req_1); -- 
    -- CP-element group 10:  transition  place  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	15 
    -- CP-element group 10:  members (7) 
      -- CP-element group 10: 	 branch_block_stmt_881/assign_stmt_960__entry__
      -- CP-element group 10: 	 branch_block_stmt_881/assign_stmt_960/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_881/assign_stmt_960/$entry
      -- CP-element group 10: 	 branch_block_stmt_881/if_stmt_945_else_link/else_choice_transition
      -- CP-element group 10: 	 branch_block_stmt_881/assign_stmt_960/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_881/assign_stmt_960/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_Sample/req
      -- CP-element group 10: 	 branch_block_stmt_881/if_stmt_945_else_link/$exit
      -- 
    else_choice_transition_1421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_945_branch_ack_0, ack => populateRxQueue_CP_1330_elements(10)); -- 
    req_1492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1330_elements(10), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_881/call_stmt_950/call_stmt_950_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_881/call_stmt_950/call_stmt_950_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_881/call_stmt_950/call_stmt_950_Sample/cra
      -- 
    cra_1437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_950_call_ack_0, ack => populateRxQueue_CP_1330_elements(11)); -- 
    -- CP-element group 12:  branch  transition  place  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (27) 
      -- CP-element group 12: 	 branch_block_stmt_881/call_stmt_950__exit__
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_eval_test/EQ_u1_u1_954/SplitProtocol/Update/ca
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_eval_test/EQ_u1_u1_954/SplitProtocol/Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_eval_test/EQ_u1_u1_954/SplitProtocol/$exit
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_eval_test/EQ_u1_u1_954/EQ_u1_u1_954_inputs/$exit
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_if_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_881/call_stmt_950/call_stmt_950_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_eval_test/EQ_u1_u1_954/SplitProtocol/Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_eval_test/branch_req
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_eval_test/EQ_u1_u1_954/SplitProtocol/Update/cr
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_eval_test/EQ_u1_u1_954/SplitProtocol/Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_eval_test/EQ_u1_u1_954/SplitProtocol/Sample/rr
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_eval_test/EQ_u1_u1_954/SplitProtocol/Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_eval_test/EQ_u1_u1_954/SplitProtocol/$entry
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_eval_test/$entry
      -- CP-element group 12: 	 branch_block_stmt_881/EQ_u1_u1_954_place
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_dead_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_else_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_eval_test/EQ_u1_u1_954/EQ_u1_u1_954_inputs/$entry
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951__entry__
      -- CP-element group 12: 	 branch_block_stmt_881/call_stmt_950/$exit
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_eval_test/EQ_u1_u1_954/$exit
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_eval_test/EQ_u1_u1_954/SplitProtocol/Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_eval_test/EQ_u1_u1_954/$entry
      -- CP-element group 12: 	 branch_block_stmt_881/if_stmt_951_eval_test/$exit
      -- CP-element group 12: 	 branch_block_stmt_881/call_stmt_950/call_stmt_950_Update/cca
      -- CP-element group 12: 	 branch_block_stmt_881/call_stmt_950/call_stmt_950_Update/$exit
      -- 
    cca_1442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_950_call_ack_1, ack => populateRxQueue_CP_1330_elements(12)); -- 
    branch_req_1469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1330_elements(12), ack => if_stmt_951_branch_req_0); -- 
    -- CP-element group 13:  fork  transition  place  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	21 
    -- CP-element group 13: 	22 
    -- CP-element group 13:  members (11) 
      -- CP-element group 13: 	 branch_block_stmt_881/loopback_PhiReq/phi_stmt_883/phi_stmt_883_sources/Interlock/$entry
      -- CP-element group 13: 	 branch_block_stmt_881/loopback_PhiReq/phi_stmt_883/phi_stmt_883_sources/Interlock/Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_881/loopback_PhiReq/phi_stmt_883/$entry
      -- CP-element group 13: 	 branch_block_stmt_881/loopback_PhiReq/$entry
      -- CP-element group 13: 	 branch_block_stmt_881/if_stmt_951_if_link/$exit
      -- CP-element group 13: 	 branch_block_stmt_881/loopback
      -- CP-element group 13: 	 branch_block_stmt_881/if_stmt_951_if_link/if_choice_transition
      -- CP-element group 13: 	 branch_block_stmt_881/loopback_PhiReq/phi_stmt_883/phi_stmt_883_sources/$entry
      -- CP-element group 13: 	 branch_block_stmt_881/loopback_PhiReq/phi_stmt_883/phi_stmt_883_sources/Interlock/Update/req
      -- CP-element group 13: 	 branch_block_stmt_881/loopback_PhiReq/phi_stmt_883/phi_stmt_883_sources/Interlock/Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_881/loopback_PhiReq/phi_stmt_883/phi_stmt_883_sources/Interlock/Sample/req
      -- 
    if_choice_transition_1474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_951_branch_ack_1, ack => populateRxQueue_CP_1330_elements(13)); -- 
    req_1632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1330_elements(13), ack => n_q_index_941_893_buf_req_1); -- 
    req_1627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1330_elements(13), ack => n_q_index_941_893_buf_req_0); -- 
    -- CP-element group 14:  merge  transition  place  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	1 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_881/if_stmt_951__exit__
      -- CP-element group 14: 	 branch_block_stmt_881/if_stmt_951_else_link/else_choice_transition
      -- CP-element group 14: 	 branch_block_stmt_881/if_stmt_951_else_link/$exit
      -- 
    else_choice_transition_1478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_951_branch_ack_0, ack => populateRxQueue_CP_1330_elements(14)); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_881/assign_stmt_960/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_update_start_
      -- CP-element group 15: 	 branch_block_stmt_881/assign_stmt_960/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_Update/req
      -- CP-element group 15: 	 branch_block_stmt_881/assign_stmt_960/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_881/assign_stmt_960/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_Sample/ack
      -- CP-element group 15: 	 branch_block_stmt_881/assign_stmt_960/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_881/assign_stmt_960/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_Update/$entry
      -- 
    ack_1493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_inst_ack_0, ack => populateRxQueue_CP_1330_elements(15)); -- 
    req_1497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1330_elements(15), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_inst_req_1); -- 
    -- CP-element group 16:  transition  place  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	1 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_881/assign_stmt_960/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_Update/ack
      -- CP-element group 16: 	 branch_block_stmt_881/assign_stmt_960/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_881/assign_stmt_960__exit__
      -- CP-element group 16: 	 branch_block_stmt_881/assign_stmt_960/$exit
      -- CP-element group 16: 	 branch_block_stmt_881/assign_stmt_960/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_Update/$exit
      -- 
    ack_1498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_inst_ack_1, ack => populateRxQueue_CP_1330_elements(16)); -- 
    -- CP-element group 17:  join  fork  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (71) 
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/SplitProtocol/Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SplitProtocol/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/SplitProtocol/Update/ca
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SUB_u32_u32_890_inputs/RPIPE_NUMBER_OF_SERVERS_888/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/SplitProtocol/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SplitProtocol/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SplitProtocol/Update/ca
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SplitProtocol/Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SUB_u32_u32_890_inputs/RPIPE_NUMBER_OF_SERVERS_888/Sample/req
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/SplitProtocol/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SUB_u32_u32_890_inputs/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/SplitProtocol/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SplitProtocol/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SUB_u32_u32_890_inputs/RPIPE_NUMBER_OF_SERVERS_888/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SplitProtocol/Update/cr
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SplitProtocol/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SplitProtocol/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/SplitProtocol/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/SplitProtocol/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SUB_u32_u32_890_inputs/RPIPE_NUMBER_OF_SERVERS_888/Update/ack
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/SplitProtocol/Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/SplitProtocol/Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SplitProtocol/Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SUB_u32_u32_890_inputs/RPIPE_NUMBER_OF_SERVERS_888/Sample/ack
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SUB_u32_u32_890_inputs/RPIPE_NUMBER_OF_SERVERS_888/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SplitProtocol/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/ADD_u6_u6_887_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_885/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/SplitProtocol/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/SplitProtocol/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SplitProtocol/Update/ca
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SplitProtocol/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SplitProtocol/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SplitProtocol/Update/cr
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SplitProtocol/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SplitProtocol/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/SplitProtocol/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SUB_u32_u32_890_inputs/RPIPE_NUMBER_OF_SERVERS_888/Update/req
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SplitProtocol/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/ADD_u6_u6_887_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_885/Update/req
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/SplitProtocol/Update/cr
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/SplitProtocol/Update/cr
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SplitProtocol/Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SplitProtocol/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/SplitProtocol/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/ADD_u6_u6_887_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_885/Update/ack
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SUB_u32_u32_890_inputs/RPIPE_NUMBER_OF_SERVERS_888/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SUB_u32_u32_890_inputs/RPIPE_NUMBER_OF_SERVERS_888/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/ADD_u6_u6_887_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_885/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/ADD_u6_u6_887_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_885/Sample/ack
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SUB_u32_u32_890_inputs/RPIPE_NUMBER_OF_SERVERS_888/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SplitProtocol/Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/ADD_u6_u6_887_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_885/Sample/req
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/ADD_u6_u6_887_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_885/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/ADD_u6_u6_887_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_885/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/ADD_u6_u6_887_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_885/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/ADD_u6_u6_887_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_885/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/ADD_u6_u6_887_inputs/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/ADD_u6_u6_887_inputs/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/ADD_u6_u6_887/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/$entry
      -- CP-element group 17: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/AND_u6_u6_892_inputs/type_cast_891/SUB_u32_u32_890/SUB_u32_u32_890_inputs/$exit
      -- 
    rr_1604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1330_elements(17), ack => AND_u6_u6_892_inst_req_0); -- 
    cr_1609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1330_elements(17), ack => AND_u6_u6_892_inst_req_1); -- 
    populateRxQueue_CP_1330_elements(17) <= populateRxQueue_CP_1330_elements(0);
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/SplitProtocol/Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/SplitProtocol/Sample/$exit
      -- 
    ra_1605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_892_inst_ack_0, ack => populateRxQueue_CP_1330_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/SplitProtocol/Update/ca
      -- CP-element group 19: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/SplitProtocol/Update/$exit
      -- 
    ca_1610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_892_inst_ack_1, ack => populateRxQueue_CP_1330_elements(19)); -- 
    -- CP-element group 20:  join  transition  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	24 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/SplitProtocol/$exit
      -- CP-element group 20: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/$exit
      -- CP-element group 20: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/$exit
      -- CP-element group 20: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_req
      -- CP-element group 20: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/$exit
      -- CP-element group 20: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/phi_stmt_883/phi_stmt_883_sources/AND_u6_u6_892/$exit
      -- 
    phi_stmt_883_req_1611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_883_req_1611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1330_elements(20), ack => phi_stmt_883_req_0); -- 
    populateRxQueue_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "populateRxQueue_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_1330_elements(18) & populateRxQueue_CP_1330_elements(19);
      gj_populateRxQueue_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_1330_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	13 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_881/loopback_PhiReq/phi_stmt_883/phi_stmt_883_sources/Interlock/Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_881/loopback_PhiReq/phi_stmt_883/phi_stmt_883_sources/Interlock/Sample/ack
      -- 
    ack_1628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_q_index_941_893_buf_ack_0, ack => populateRxQueue_CP_1330_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	13 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_881/loopback_PhiReq/phi_stmt_883/phi_stmt_883_sources/Interlock/Update/ack
      -- CP-element group 22: 	 branch_block_stmt_881/loopback_PhiReq/phi_stmt_883/phi_stmt_883_sources/Interlock/Update/$exit
      -- 
    ack_1633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_q_index_941_893_buf_ack_1, ack => populateRxQueue_CP_1330_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_881/loopback_PhiReq/phi_stmt_883/phi_stmt_883_sources/$exit
      -- CP-element group 23: 	 branch_block_stmt_881/loopback_PhiReq/phi_stmt_883/$exit
      -- CP-element group 23: 	 branch_block_stmt_881/loopback_PhiReq/phi_stmt_883/phi_stmt_883_req
      -- CP-element group 23: 	 branch_block_stmt_881/loopback_PhiReq/phi_stmt_883/phi_stmt_883_sources/Interlock/$exit
      -- CP-element group 23: 	 branch_block_stmt_881/loopback_PhiReq/$exit
      -- 
    phi_stmt_883_req_1634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_883_req_1634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1330_elements(23), ack => phi_stmt_883_req_1); -- 
    populateRxQueue_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "populateRxQueue_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_1330_elements(21) & populateRxQueue_CP_1330_elements(22);
      gj_populateRxQueue_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_1330_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  merge  transition  place  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	20 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_881/merge_stmt_882_PhiReqMerge
      -- CP-element group 24: 	 branch_block_stmt_881/merge_stmt_882_PhiAck/$entry
      -- 
    populateRxQueue_CP_1330_elements(24) <= OrReduce(populateRxQueue_CP_1330_elements(20) & populateRxQueue_CP_1330_elements(23));
    -- CP-element group 25:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: 	3 
    -- CP-element group 25: 	5 
    -- CP-element group 25: 	6 
    -- CP-element group 25: 	7 
    -- CP-element group 25:  members (20) 
      -- CP-element group 25: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_931_Update/ccr
      -- CP-element group 25: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_914_Sample/crr
      -- CP-element group 25: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_931_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_914_update_start_
      -- CP-element group 25: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_914_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941__entry__
      -- CP-element group 25: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/$entry
      -- CP-element group 25: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/AND_u6_u6_940_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_931_update_start_
      -- CP-element group 25: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_914_Update/ccr
      -- CP-element group 25: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_914_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/call_stmt_914_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/AND_u6_u6_940_Update/cr
      -- CP-element group 25: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/AND_u6_u6_940_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_881/merge_stmt_882_PhiAck/phi_stmt_883_ack
      -- CP-element group 25: 	 branch_block_stmt_881/merge_stmt_882_PhiAck/$exit
      -- CP-element group 25: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/AND_u6_u6_940_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/AND_u6_u6_940_update_start_
      -- CP-element group 25: 	 branch_block_stmt_881/assign_stmt_902_to_assign_stmt_941/AND_u6_u6_940_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_881/merge_stmt_882__exit__
      -- 
    phi_stmt_883_ack_1639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_883_ack_0, ack => populateRxQueue_CP_1330_elements(25)); -- 
    ccr_1373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1330_elements(25), ack => call_stmt_931_call_req_1); -- 
    crr_1354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1330_elements(25), ack => call_stmt_914_call_req_0); -- 
    ccr_1359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1330_elements(25), ack => call_stmt_914_call_req_1); -- 
    cr_1387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1330_elements(25), ack => AND_u6_u6_940_inst_req_1); -- 
    rr_1382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1330_elements(25), ack => AND_u6_u6_940_inst_req_0); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u6_u6_887_wire : std_logic_vector(5 downto 0);
    signal ADD_u6_u6_900_wire : std_logic_vector(5 downto 0);
    signal ADD_u6_u6_935_wire : std_logic_vector(5 downto 0);
    signal AND_u6_u6_892_wire : std_logic_vector(5 downto 0);
    signal EQ_u1_u1_954_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_947_wire : std_logic_vector(0 downto 0);
    signal NOT_u4_u4_909_wire_constant : std_logic_vector(3 downto 0);
    signal RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_885_wire : std_logic_vector(5 downto 0);
    signal RPIPE_NUMBER_OF_SERVERS_888_wire : std_logic_vector(31 downto 0);
    signal RPIPE_NUMBER_OF_SERVERS_936_wire : std_logic_vector(31 downto 0);
    signal R_RX_QUEUES_REG_START_OFFSET_899_wire_constant : std_logic_vector(5 downto 0);
    signal SUB_u32_u32_890_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_938_wire : std_logic_vector(31 downto 0);
    signal konst_886_wire_constant : std_logic_vector(5 downto 0);
    signal konst_889_wire_constant : std_logic_vector(31 downto 0);
    signal konst_934_wire_constant : std_logic_vector(5 downto 0);
    signal konst_937_wire_constant : std_logic_vector(31 downto 0);
    signal konst_948_wire_constant : std_logic_vector(31 downto 0);
    signal konst_953_wire_constant : std_logic_vector(0 downto 0);
    signal n_q_index_941 : std_logic_vector(5 downto 0);
    signal n_q_index_941_893_buffered : std_logic_vector(5 downto 0);
    signal push_status_931 : std_logic_vector(0 downto 0);
    signal q_index_883 : std_logic_vector(5 downto 0);
    signal register_index_902 : std_logic_vector(5 downto 0);
    signal rx_queue_pointer_32_914 : std_logic_vector(31 downto 0);
    signal rx_queue_pointer_36_920 : std_logic_vector(35 downto 0);
    signal slice_929_wire : std_logic_vector(31 downto 0);
    signal status_950 : std_logic_vector(0 downto 0);
    signal type_cast_891_wire : std_logic_vector(5 downto 0);
    signal type_cast_906_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_912_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_918_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_926_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_939_wire : std_logic_vector(5 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_909_wire_constant <= "1111";
    R_RX_QUEUES_REG_START_OFFSET_899_wire_constant <= "000010";
    konst_886_wire_constant <= "000001";
    konst_889_wire_constant <= "00000000000000000000000000000001";
    konst_934_wire_constant <= "000001";
    konst_937_wire_constant <= "00000000000000000000000000000001";
    konst_948_wire_constant <= "00000000000000000000000000100000";
    konst_953_wire_constant <= "0";
    type_cast_906_wire_constant <= "1";
    type_cast_912_wire_constant <= "00000000000000000000000000000000";
    type_cast_918_wire_constant <= "0000";
    type_cast_926_wire_constant <= "0";
    phi_stmt_883: Block -- phi operator 
      signal idata: std_logic_vector(11 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= AND_u6_u6_892_wire & n_q_index_941_893_buffered;
      req <= phi_stmt_883_req_0 & phi_stmt_883_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_883",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 6) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_883_ack_0,
          idata => idata,
          odata => q_index_883,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_883
    -- flow-through slice operator slice_929_inst
    slice_929_wire <= rx_buffer_pointer_buffer(35 downto 4);
    n_q_index_941_893_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_q_index_941_893_buf_req_0;
      n_q_index_941_893_buf_ack_0<= wack(0);
      rreq(0) <= n_q_index_941_893_buf_req_1;
      n_q_index_941_893_buf_ack_1<= rack(0);
      n_q_index_941_893_buf : InterlockBuffer generic map ( -- 
        name => "n_q_index_941_893_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_q_index_941,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_q_index_941_893_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_891_inst
    process(SUB_u32_u32_890_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := SUB_u32_u32_890_wire(5 downto 0);
      type_cast_891_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_901_inst
    process(ADD_u6_u6_900_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := ADD_u6_u6_900_wire(5 downto 0);
      register_index_902 <= tmp_var; -- 
    end process;
    -- interlock type_cast_939_inst
    process(SUB_u32_u32_938_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := SUB_u32_u32_938_wire(5 downto 0);
      type_cast_939_wire <= tmp_var; -- 
    end process;
    if_stmt_945_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_947_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_945_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_945_branch_req_0,
          ack0 => if_stmt_945_branch_ack_0,
          ack1 => if_stmt_945_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_951_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_954_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_951_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_951_branch_req_0,
          ack0 => if_stmt_951_branch_ack_0,
          ack1 => if_stmt_951_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u6_u6_887_inst
    process(RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_885_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_885_wire, konst_886_wire_constant, tmp_var);
      ADD_u6_u6_887_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u6_u6_900_inst
    process(q_index_883) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_index_883, R_RX_QUEUES_REG_START_OFFSET_899_wire_constant, tmp_var);
      ADD_u6_u6_900_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u6_u6_935_inst
    process(q_index_883) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_index_883, konst_934_wire_constant, tmp_var);
      ADD_u6_u6_935_wire <= tmp_var; --
    end process;
    -- shared split operator group (3) : AND_u6_u6_892_inst 
    ApIntAnd_group_3: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u6_u6_887_wire & type_cast_891_wire;
      AND_u6_u6_892_wire <= data_out(5 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u6_u6_892_inst_req_0;
      AND_u6_u6_892_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u6_u6_892_inst_req_1;
      AND_u6_u6_892_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 6, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : AND_u6_u6_940_inst 
    ApIntAnd_group_4: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u6_u6_935_wire & type_cast_939_wire;
      n_q_index_941 <= data_out(5 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u6_u6_940_inst_req_0;
      AND_u6_u6_940_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u6_u6_940_inst_req_1;
      AND_u6_u6_940_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_4_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 6, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- binary operator CONCAT_u32_u36_919_inst
    process(rx_queue_pointer_32_914) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(rx_queue_pointer_32_914, type_cast_918_wire_constant, tmp_var);
      rx_queue_pointer_36_920 <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_954_inst
    process(status_950) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(status_950, konst_953_wire_constant, tmp_var);
      EQ_u1_u1_954_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_947_inst
    process(push_status_931) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", push_status_931, tmp_var);
      NOT_u1_u1_947_wire <= tmp_var; -- 
    end process;
    -- binary operator SUB_u32_u32_890_inst
    process(RPIPE_NUMBER_OF_SERVERS_888_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(RPIPE_NUMBER_OF_SERVERS_888_wire, konst_889_wire_constant, tmp_var);
      SUB_u32_u32_890_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_938_inst
    process(RPIPE_NUMBER_OF_SERVERS_936_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(RPIPE_NUMBER_OF_SERVERS_936_wire, konst_937_wire_constant, tmp_var);
      SUB_u32_u32_938_wire <= tmp_var; --
    end process;
    -- read from input-signal LAST_WRITTEN_RX_QUEUE_INDEX
    RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_885_wire <= LAST_WRITTEN_RX_QUEUE_INDEX;
    -- read from input-signal NUMBER_OF_SERVERS
    RPIPE_NUMBER_OF_SERVERS_888_wire <= NUMBER_OF_SERVERS;
    RPIPE_NUMBER_OF_SERVERS_936_wire <= NUMBER_OF_SERVERS;
    -- shared outport operator group (0) : WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_inst_req_0;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_inst_req_1;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_958_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= q_index_883;
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_WRITTEN_RX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(5 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_914_call 
    AccessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_914_call_req_0;
      call_stmt_914_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_914_call_req_1;
      call_stmt_914_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_906_wire_constant & NOT_u4_u4_909_wire_constant & register_index_902 & type_cast_912_wire_constant;
      rx_queue_pointer_32_914 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_931_call 
    pushIntoQueue_call_group_1: Block -- 
      signal data_in: std_logic_vector(68 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_931_call_req_0;
      call_stmt_931_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_931_call_req_1;
      call_stmt_931_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_1_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_926_wire_constant & rx_queue_pointer_36_920 & slice_929_wire;
      push_status_931 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 69,
        owidth => 69,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(68 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    operator_delay_time_2323_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_950_call_req_0;
      call_stmt_950_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_950_call_req_1;
      call_stmt_950_call_ack_1<= update_ack(0);
      call_stmt_950_call: delay_time_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        T => konst_948_wire_constant,
        delay_done => status_950,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- 
  end Block; -- data_path
  -- 
end populateRxQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity pushIntoQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    lock : in  std_logic_vector(0 downto 0);
    q_base_address : in  std_logic_vector(35 downto 0);
    q_w_data : in  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
    setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
    releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
    releaseMutex_call_data : out  std_logic_vector(35 downto 0);
    releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
    releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
    releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
    releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
    getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
    getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
    getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
    acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
    acquireMutex_call_data : out  std_logic_vector(35 downto 0);
    acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
    acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
    acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
    acquireMutex_return_data : in   std_logic_vector(0 downto 0);
    acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
    setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
    setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
    setQueueElement_call_data : out  std_logic_vector(99 downto 0);
    setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
    setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
    setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity pushIntoQueue;
architecture pushIntoQueue_arch of pushIntoQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 69)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal q_w_data_buffer :  std_logic_vector(31 downto 0);
  signal q_w_data_update_enable: Boolean;
  -- output port buffer signals
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal pushIntoQueue_CP_1135_start: Boolean;
  signal pushIntoQueue_CP_1135_symbol: Boolean;
  -- volatile/operator module components. 
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component releaseMutex is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component acquireMutex is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component setQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      write_pointer : in  std_logic_vector(31 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_798_call_req_0 : boolean;
  signal call_stmt_798_call_ack_0 : boolean;
  signal call_stmt_798_call_req_1 : boolean;
  signal call_stmt_798_call_ack_1 : boolean;
  signal call_stmt_806_call_req_0 : boolean;
  signal call_stmt_806_call_ack_0 : boolean;
  signal call_stmt_806_call_req_1 : boolean;
  signal call_stmt_806_call_ack_1 : boolean;
  signal call_stmt_837_call_req_0 : boolean;
  signal call_stmt_837_call_ack_0 : boolean;
  signal call_stmt_837_call_req_1 : boolean;
  signal call_stmt_837_call_ack_1 : boolean;
  signal call_stmt_842_call_req_0 : boolean;
  signal call_stmt_842_call_ack_0 : boolean;
  signal call_stmt_842_call_req_1 : boolean;
  signal call_stmt_842_call_ack_1 : boolean;
  signal call_stmt_846_call_req_0 : boolean;
  signal call_stmt_846_call_ack_0 : boolean;
  signal call_stmt_846_call_req_1 : boolean;
  signal call_stmt_846_call_ack_1 : boolean;
  signal NOT_u1_u1_849_inst_req_0 : boolean;
  signal NOT_u1_u1_849_inst_ack_0 : boolean;
  signal NOT_u1_u1_849_inst_req_1 : boolean;
  signal NOT_u1_u1_849_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "pushIntoQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 69) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= lock;
  lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(36 downto 1) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(36 downto 1);
  in_buffer_data_in(68 downto 37) <= q_w_data;
  q_w_data_buffer <= in_buffer_data_out(68 downto 37);
  in_buffer_data_in(tag_length + 68 downto 69) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 68 downto 69);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  pushIntoQueue_CP_1135_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "pushIntoQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= status_buffer;
  status <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= pushIntoQueue_CP_1135_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= pushIntoQueue_CP_1135_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= pushIntoQueue_CP_1135_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  pushIntoQueue_CP_1135: Block -- control-path 
    signal pushIntoQueue_CP_1135_elements: BooleanArray(14 downto 0);
    -- 
  begin -- 
    pushIntoQueue_CP_1135_elements(0) <= pushIntoQueue_CP_1135_start;
    pushIntoQueue_CP_1135_symbol <= pushIntoQueue_CP_1135_elements(14);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_798/$entry
      -- CP-element group 0: 	 call_stmt_798/call_stmt_798_sample_start_
      -- CP-element group 0: 	 call_stmt_798/call_stmt_798_update_start_
      -- CP-element group 0: 	 call_stmt_798/call_stmt_798_Sample/$entry
      -- CP-element group 0: 	 call_stmt_798/call_stmt_798_Sample/crr
      -- CP-element group 0: 	 call_stmt_798/call_stmt_798_Update/$entry
      -- CP-element group 0: 	 call_stmt_798/call_stmt_798_Update/ccr
      -- 
    crr_1148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1135_elements(0), ack => call_stmt_798_call_req_0); -- 
    ccr_1153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1135_elements(0), ack => call_stmt_798_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_798/call_stmt_798_sample_completed_
      -- CP-element group 1: 	 call_stmt_798/call_stmt_798_Sample/$exit
      -- CP-element group 1: 	 call_stmt_798/call_stmt_798_Sample/cra
      -- 
    cra_1149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_798_call_ack_0, ack => pushIntoQueue_CP_1135_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	9 
    -- CP-element group 2:  members (17) 
      -- CP-element group 2: 	 call_stmt_798/$exit
      -- CP-element group 2: 	 call_stmt_798/call_stmt_798_update_completed_
      -- CP-element group 2: 	 call_stmt_798/call_stmt_798_Update/$exit
      -- CP-element group 2: 	 call_stmt_798/call_stmt_798_Update/cca
      -- CP-element group 2: 	 call_stmt_806_to_call_stmt_842/$entry
      -- CP-element group 2: 	 call_stmt_806_to_call_stmt_842/call_stmt_806_sample_start_
      -- CP-element group 2: 	 call_stmt_806_to_call_stmt_842/call_stmt_806_update_start_
      -- CP-element group 2: 	 call_stmt_806_to_call_stmt_842/call_stmt_806_Sample/$entry
      -- CP-element group 2: 	 call_stmt_806_to_call_stmt_842/call_stmt_806_Sample/crr
      -- CP-element group 2: 	 call_stmt_806_to_call_stmt_842/call_stmt_806_Update/$entry
      -- CP-element group 2: 	 call_stmt_806_to_call_stmt_842/call_stmt_806_Update/ccr
      -- CP-element group 2: 	 call_stmt_806_to_call_stmt_842/call_stmt_837_update_start_
      -- CP-element group 2: 	 call_stmt_806_to_call_stmt_842/call_stmt_837_Update/$entry
      -- CP-element group 2: 	 call_stmt_806_to_call_stmt_842/call_stmt_837_Update/ccr
      -- CP-element group 2: 	 call_stmt_806_to_call_stmt_842/call_stmt_842_update_start_
      -- CP-element group 2: 	 call_stmt_806_to_call_stmt_842/call_stmt_842_Update/$entry
      -- CP-element group 2: 	 call_stmt_806_to_call_stmt_842/call_stmt_842_Update/ccr
      -- 
    cca_1154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_798_call_ack_1, ack => pushIntoQueue_CP_1135_elements(2)); -- 
    crr_1165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1135_elements(2), ack => call_stmt_806_call_req_0); -- 
    ccr_1170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1135_elements(2), ack => call_stmt_806_call_req_1); -- 
    ccr_1184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1135_elements(2), ack => call_stmt_837_call_req_1); -- 
    ccr_1198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1135_elements(2), ack => call_stmt_842_call_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_806_to_call_stmt_842/call_stmt_806_sample_completed_
      -- CP-element group 3: 	 call_stmt_806_to_call_stmt_842/call_stmt_806_Sample/$exit
      -- CP-element group 3: 	 call_stmt_806_to_call_stmt_842/call_stmt_806_Sample/cra
      -- 
    cra_1166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_806_call_ack_0, ack => pushIntoQueue_CP_1135_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 call_stmt_806_to_call_stmt_842/call_stmt_806_update_completed_
      -- CP-element group 4: 	 call_stmt_806_to_call_stmt_842/call_stmt_806_Update/$exit
      -- CP-element group 4: 	 call_stmt_806_to_call_stmt_842/call_stmt_806_Update/cca
      -- CP-element group 4: 	 call_stmt_806_to_call_stmt_842/call_stmt_837_sample_start_
      -- CP-element group 4: 	 call_stmt_806_to_call_stmt_842/call_stmt_837_Sample/$entry
      -- CP-element group 4: 	 call_stmt_806_to_call_stmt_842/call_stmt_837_Sample/crr
      -- 
    cca_1171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_806_call_ack_1, ack => pushIntoQueue_CP_1135_elements(4)); -- 
    crr_1179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1135_elements(4), ack => call_stmt_837_call_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_806_to_call_stmt_842/call_stmt_837_sample_completed_
      -- CP-element group 5: 	 call_stmt_806_to_call_stmt_842/call_stmt_837_Sample/$exit
      -- CP-element group 5: 	 call_stmt_806_to_call_stmt_842/call_stmt_837_Sample/cra
      -- 
    cra_1180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_837_call_ack_0, ack => pushIntoQueue_CP_1135_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 call_stmt_806_to_call_stmt_842/call_stmt_837_update_completed_
      -- CP-element group 6: 	 call_stmt_806_to_call_stmt_842/call_stmt_837_Update/$exit
      -- CP-element group 6: 	 call_stmt_806_to_call_stmt_842/call_stmt_837_Update/cca
      -- 
    cca_1185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_837_call_ack_1, ack => pushIntoQueue_CP_1135_elements(6)); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_806_to_call_stmt_842/call_stmt_842_sample_start_
      -- CP-element group 7: 	 call_stmt_806_to_call_stmt_842/call_stmt_842_Sample/$entry
      -- CP-element group 7: 	 call_stmt_806_to_call_stmt_842/call_stmt_842_Sample/crr
      -- 
    crr_1193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1135_elements(7), ack => call_stmt_842_call_req_0); -- 
    pushIntoQueue_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "pushIntoQueue_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= pushIntoQueue_CP_1135_elements(4) & pushIntoQueue_CP_1135_elements(6);
      gj_pushIntoQueue_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_1135_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_806_to_call_stmt_842/call_stmt_842_sample_completed_
      -- CP-element group 8: 	 call_stmt_806_to_call_stmt_842/call_stmt_842_Sample/$exit
      -- CP-element group 8: 	 call_stmt_806_to_call_stmt_842/call_stmt_842_Sample/cra
      -- 
    cra_1194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_842_call_ack_0, ack => pushIntoQueue_CP_1135_elements(8)); -- 
    -- CP-element group 9:  fork  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9:  members (17) 
      -- CP-element group 9: 	 call_stmt_806_to_call_stmt_842/$exit
      -- CP-element group 9: 	 call_stmt_806_to_call_stmt_842/call_stmt_842_update_completed_
      -- CP-element group 9: 	 call_stmt_806_to_call_stmt_842/call_stmt_842_Update/$exit
      -- CP-element group 9: 	 call_stmt_806_to_call_stmt_842/call_stmt_842_Update/cca
      -- CP-element group 9: 	 call_stmt_846_to_assign_stmt_850/$entry
      -- CP-element group 9: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_sample_start_
      -- CP-element group 9: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_update_start_
      -- CP-element group 9: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_Sample/$entry
      -- CP-element group 9: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_Sample/crr
      -- CP-element group 9: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_Update/$entry
      -- CP-element group 9: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_Update/ccr
      -- CP-element group 9: 	 call_stmt_846_to_assign_stmt_850/NOT_u1_u1_849_sample_start_
      -- CP-element group 9: 	 call_stmt_846_to_assign_stmt_850/NOT_u1_u1_849_update_start_
      -- CP-element group 9: 	 call_stmt_846_to_assign_stmt_850/NOT_u1_u1_849_Sample/$entry
      -- CP-element group 9: 	 call_stmt_846_to_assign_stmt_850/NOT_u1_u1_849_Sample/rr
      -- CP-element group 9: 	 call_stmt_846_to_assign_stmt_850/NOT_u1_u1_849_Update/$entry
      -- CP-element group 9: 	 call_stmt_846_to_assign_stmt_850/NOT_u1_u1_849_Update/cr
      -- 
    cca_1199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_842_call_ack_1, ack => pushIntoQueue_CP_1135_elements(9)); -- 
    crr_1210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1135_elements(9), ack => call_stmt_846_call_req_0); -- 
    ccr_1215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1135_elements(9), ack => call_stmt_846_call_req_1); -- 
    rr_1224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1135_elements(9), ack => NOT_u1_u1_849_inst_req_0); -- 
    cr_1229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1135_elements(9), ack => NOT_u1_u1_849_inst_req_1); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_sample_completed_
      -- CP-element group 10: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_Sample/$exit
      -- CP-element group 10: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_Sample/cra
      -- 
    cra_1211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_846_call_ack_0, ack => pushIntoQueue_CP_1135_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_update_completed_
      -- CP-element group 11: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_Update/$exit
      -- CP-element group 11: 	 call_stmt_846_to_assign_stmt_850/call_stmt_846_Update/cca
      -- 
    cca_1216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_846_call_ack_1, ack => pushIntoQueue_CP_1135_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_846_to_assign_stmt_850/NOT_u1_u1_849_sample_completed_
      -- CP-element group 12: 	 call_stmt_846_to_assign_stmt_850/NOT_u1_u1_849_Sample/$exit
      -- CP-element group 12: 	 call_stmt_846_to_assign_stmt_850/NOT_u1_u1_849_Sample/ra
      -- 
    ra_1225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_849_inst_ack_0, ack => pushIntoQueue_CP_1135_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_846_to_assign_stmt_850/NOT_u1_u1_849_update_completed_
      -- CP-element group 13: 	 call_stmt_846_to_assign_stmt_850/NOT_u1_u1_849_Update/$exit
      -- CP-element group 13: 	 call_stmt_846_to_assign_stmt_850/NOT_u1_u1_849_Update/ca
      -- 
    ca_1230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_849_inst_ack_1, ack => pushIntoQueue_CP_1135_elements(13)); -- 
    -- CP-element group 14:  join  transition  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 $exit
      -- CP-element group 14: 	 call_stmt_846_to_assign_stmt_850/$exit
      -- 
    pushIntoQueue_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= pushIntoQueue_CP_1135_elements(11) & pushIntoQueue_CP_1135_elements(13);
      gj_pushIntoQueue_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_1135_elements(14), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_819_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_811_wire_constant : std_logic_vector(31 downto 0);
    signal konst_816_wire_constant : std_logic_vector(31 downto 0);
    signal konst_818_wire_constant : std_logic_vector(31 downto 0);
    signal m_ok_798 : std_logic_vector(0 downto 0);
    signal next_wp_821 : std_logic_vector(31 downto 0);
    signal q_full_826 : std_logic_vector(0 downto 0);
    signal read_pointer_806 : std_logic_vector(31 downto 0);
    signal round_off_813 : std_logic_vector(0 downto 0);
    signal write_pointer_806 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    SUB_u32_u32_811_wire_constant <= "00000000000000000000000000000111";
    konst_816_wire_constant <= "00000000000000000000000000000000";
    konst_818_wire_constant <= "00000000000000000000000000000001";
    -- flow-through select operator MUX_820_inst
    next_wp_821 <= konst_816_wire_constant when (round_off_813(0) /=  '0') else ADD_u32_u32_819_wire;
    -- binary operator ADD_u32_u32_819_inst
    process(write_pointer_806) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(write_pointer_806, konst_818_wire_constant, tmp_var);
      ADD_u32_u32_819_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_812_inst
    process(write_pointer_806) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(write_pointer_806, SUB_u32_u32_811_wire_constant, tmp_var);
      round_off_813 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_825_inst
    process(next_wp_821, read_pointer_806) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_wp_821, read_pointer_806, tmp_var);
      q_full_826 <= tmp_var; --
    end process;
    -- shared split operator group (3) : NOT_u1_u1_849_inst 
    ApIntNot_group_3: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= q_full_826;
      status_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_849_inst_req_0;
      NOT_u1_u1_849_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_849_inst_req_1;
      NOT_u1_u1_849_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_3_gI: SplitGuardInterface generic map(name => "ApIntNot_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared call operator group (0) : call_stmt_798_call 
    acquireMutex_call_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_798_call_req_0;
      call_stmt_798_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_798_call_req_1;
      call_stmt_798_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      acquireMutex_call_group_0_gI: SplitGuardInterface generic map(name => "acquireMutex_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      m_ok_798 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => acquireMutex_call_reqs(0),
          ackR => acquireMutex_call_acks(0),
          dataR => acquireMutex_call_data(35 downto 0),
          tagR => acquireMutex_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => acquireMutex_return_acks(0), -- cross-over
          ackL => acquireMutex_return_reqs(0), -- cross-over
          dataL => acquireMutex_return_data(0 downto 0),
          tagL => acquireMutex_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_806_call 
    getQueuePointers_call_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_806_call_req_0;
      call_stmt_806_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_806_call_req_1;
      call_stmt_806_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueuePointers_call_group_1_gI: SplitGuardInterface generic map(name => "getQueuePointers_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      write_pointer_806 <= data_out(63 downto 32);
      read_pointer_806 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueuePointers_call_reqs(0),
          ackR => getQueuePointers_call_acks(0),
          dataR => getQueuePointers_call_data(35 downto 0),
          tagR => getQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueuePointers_return_acks(0), -- cross-over
          ackL => getQueuePointers_return_reqs(0), -- cross-over
          dataL => getQueuePointers_return_data(63 downto 0),
          tagL => getQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_837_call 
    setQueueElement_call_group_2: Block -- 
      signal data_in: std_logic_vector(99 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_837_call_req_0;
      call_stmt_837_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_837_call_req_1;
      call_stmt_837_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_826(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueueElement_call_group_2_gI: SplitGuardInterface generic map(name => "setQueueElement_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & write_pointer_806 & q_w_data_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 100,
        owidth => 100,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueueElement_call_reqs(0),
          ackR => setQueueElement_call_acks(0),
          dataR => setQueueElement_call_data(99 downto 0),
          tagR => setQueueElement_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueueElement_return_acks(0), -- cross-over
          ackL => setQueueElement_return_reqs(0), -- cross-over
          tagL => setQueueElement_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_842_call 
    setQueuePointers_call_group_3: Block -- 
      signal data_in: std_logic_vector(99 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_842_call_req_0;
      call_stmt_842_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_842_call_req_1;
      call_stmt_842_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_826(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueuePointers_call_group_3_gI: SplitGuardInterface generic map(name => "setQueuePointers_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & next_wp_821 & read_pointer_806;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 100,
        owidth => 100,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueuePointers_call_reqs(0),
          ackR => setQueuePointers_call_acks(0),
          dataR => setQueuePointers_call_data(99 downto 0),
          tagR => setQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueuePointers_return_acks(0), -- cross-over
          ackL => setQueuePointers_return_reqs(0), -- cross-over
          tagL => setQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_846_call 
    releaseMutex_call_group_4: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_846_call_req_0;
      call_stmt_846_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_846_call_req_1;
      call_stmt_846_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      releaseMutex_call_group_4_gI: SplitGuardInterface generic map(name => "releaseMutex_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => releaseMutex_call_reqs(0),
          ackR => releaseMutex_call_acks(0),
          dataR => releaseMutex_call_data(35 downto 0),
          tagR => releaseMutex_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => releaseMutex_return_acks(0), -- cross-over
          ackL => releaseMutex_return_reqs(0), -- cross-over
          tagL => releaseMutex_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- 
  end Block; -- data_path
  -- 
end pushIntoQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity releaseMutex is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity releaseMutex;
architecture releaseMutex_arch of releaseMutex is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal releaseMutex_CP_584_start: Boolean;
  signal releaseMutex_CP_584_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_482_call_req_0 : boolean;
  signal call_stmt_482_call_ack_0 : boolean;
  signal call_stmt_482_call_req_1 : boolean;
  signal call_stmt_482_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "releaseMutex_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  releaseMutex_CP_584_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "releaseMutex_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= releaseMutex_CP_584_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= releaseMutex_CP_584_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= releaseMutex_CP_584_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  releaseMutex_CP_584: Block -- control-path 
    signal releaseMutex_CP_584_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    releaseMutex_CP_584_elements(0) <= releaseMutex_CP_584_start;
    releaseMutex_CP_584_symbol <= releaseMutex_CP_584_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_482/call_stmt_482_Sample/crr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_482/call_stmt_482_Update/$entry
      -- CP-element group 0: 	 call_stmt_482/call_stmt_482_Sample/$entry
      -- CP-element group 0: 	 call_stmt_482/call_stmt_482_Update/ccr
      -- CP-element group 0: 	 call_stmt_482/call_stmt_482_update_start_
      -- CP-element group 0: 	 call_stmt_482/$entry
      -- CP-element group 0: 	 call_stmt_482/call_stmt_482_sample_start_
      -- 
    crr_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseMutex_CP_584_elements(0), ack => call_stmt_482_call_req_0); -- 
    ccr_602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseMutex_CP_584_elements(0), ack => call_stmt_482_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_482/call_stmt_482_Sample/cra
      -- CP-element group 1: 	 call_stmt_482/call_stmt_482_Sample/$exit
      -- CP-element group 1: 	 call_stmt_482/call_stmt_482_sample_completed_
      -- 
    cra_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_482_call_ack_0, ack => releaseMutex_CP_584_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_482/$exit
      -- CP-element group 2: 	 call_stmt_482/call_stmt_482_Update/$exit
      -- CP-element group 2: 	 call_stmt_482/call_stmt_482_Update/cca
      -- CP-element group 2: 	 call_stmt_482/call_stmt_482_update_completed_
      -- 
    cca_603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_482_call_ack_1, ack => releaseMutex_CP_584_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u4_u8_477_wire_constant : std_logic_vector(7 downto 0);
    signal ignore_482 : std_logic_vector(63 downto 0);
    signal type_cast_469_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_471_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_480_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    CONCAT_u4_u8_477_wire_constant <= "11110000";
    type_cast_469_wire_constant <= "0";
    type_cast_471_wire_constant <= "0";
    type_cast_480_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- shared call operator group (0) : call_stmt_482_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_482_call_req_0;
      call_stmt_482_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_482_call_req_1;
      call_stmt_482_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_469_wire_constant & type_cast_471_wire_constant & CONCAT_u4_u8_477_wire_constant & q_base_address_buffer & type_cast_480_wire_constant;
      ignore_482 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end releaseMutex_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity setQueueElement is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    write_pointer : in  std_logic_vector(31 downto 0);
    q_w_data : in  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity setQueueElement;
architecture setQueueElement_arch of setQueueElement is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 100)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal write_pointer_buffer :  std_logic_vector(31 downto 0);
  signal write_pointer_update_enable: Boolean;
  signal q_w_data_buffer :  std_logic_vector(31 downto 0);
  signal q_w_data_update_enable: Boolean;
  -- output port buffer signals
  signal setQueueElement_CP_1115_start: Boolean;
  signal setQueueElement_CP_1115_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_788_call_req_0 : boolean;
  signal call_stmt_788_call_ack_0 : boolean;
  signal call_stmt_788_call_req_1 : boolean;
  signal call_stmt_788_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "setQueueElement_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 100) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= write_pointer;
  write_pointer_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(99 downto 68) <= q_w_data;
  q_w_data_buffer <= in_buffer_data_out(99 downto 68);
  in_buffer_data_in(tag_length + 99 downto 100) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 99 downto 100);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  setQueueElement_CP_1115_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "setQueueElement_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueueElement_CP_1115_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= setQueueElement_CP_1115_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueueElement_CP_1115_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  setQueueElement_CP_1115: Block -- control-path 
    signal setQueueElement_CP_1115_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    setQueueElement_CP_1115_elements(0) <= setQueueElement_CP_1115_start;
    setQueueElement_CP_1115_symbol <= setQueueElement_CP_1115_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_732_to_call_stmt_788/$entry
      -- CP-element group 0: 	 assign_stmt_732_to_call_stmt_788/call_stmt_788_sample_start_
      -- CP-element group 0: 	 assign_stmt_732_to_call_stmt_788/call_stmt_788_update_start_
      -- CP-element group 0: 	 assign_stmt_732_to_call_stmt_788/call_stmt_788_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_732_to_call_stmt_788/call_stmt_788_Sample/crr
      -- CP-element group 0: 	 assign_stmt_732_to_call_stmt_788/call_stmt_788_Update/$entry
      -- CP-element group 0: 	 assign_stmt_732_to_call_stmt_788/call_stmt_788_Update/ccr
      -- 
    crr_1128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueueElement_CP_1115_elements(0), ack => call_stmt_788_call_req_0); -- 
    ccr_1133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueueElement_CP_1115_elements(0), ack => call_stmt_788_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_732_to_call_stmt_788/call_stmt_788_sample_completed_
      -- CP-element group 1: 	 assign_stmt_732_to_call_stmt_788/call_stmt_788_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_732_to_call_stmt_788/call_stmt_788_Sample/cra
      -- 
    cra_1129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_788_call_ack_0, ack => setQueueElement_CP_1115_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_732_to_call_stmt_788/$exit
      -- CP-element group 2: 	 assign_stmt_732_to_call_stmt_788/call_stmt_788_update_completed_
      -- CP-element group 2: 	 assign_stmt_732_to_call_stmt_788/call_stmt_788_Update/$exit
      -- CP-element group 2: 	 assign_stmt_732_to_call_stmt_788/call_stmt_788_Update/cca
      -- 
    cca_1134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_788_call_ack_1, ack => setQueueElement_CP_1115_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_746_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_764_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u31_u34_739_wire : std_logic_vector(33 downto 0);
    signal CONCAT_u32_u64_768_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_772_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u4_u8_752_wire_constant : std_logic_vector(7 downto 0);
    signal CONCAT_u4_u8_758_wire_constant : std_logic_vector(7 downto 0);
    signal bmask_760 : std_logic_vector(7 downto 0);
    signal buffer_address_732 : std_logic_vector(35 downto 0);
    signal element_pair_address_742 : std_logic_vector(35 downto 0);
    signal ignore_788 : std_logic_vector(63 downto 0);
    signal konst_745_wire_constant : std_logic_vector(31 downto 0);
    signal konst_763_wire_constant : std_logic_vector(31 downto 0);
    signal slice_736_wire : std_logic_vector(30 downto 0);
    signal type_cast_730_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_738_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_740_wire : std_logic_vector(35 downto 0);
    signal type_cast_766_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_771_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_781_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_783_wire_constant : std_logic_vector(0 downto 0);
    signal wval_774 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    CONCAT_u4_u8_752_wire_constant <= "00001111";
    CONCAT_u4_u8_758_wire_constant <= "11110000";
    konst_745_wire_constant <= "00000000000000000000000000000000";
    konst_763_wire_constant <= "00000000000000000000000000000000";
    type_cast_730_wire_constant <= "000000000000000000000000000000010000";
    type_cast_738_wire_constant <= "000";
    type_cast_766_wire_constant <= "00000000000000000000000000000000";
    type_cast_771_wire_constant <= "00000000000000000000000000000000";
    type_cast_781_wire_constant <= "0";
    type_cast_783_wire_constant <= "0";
    -- flow-through select operator MUX_759_inst
    bmask_760 <= CONCAT_u4_u8_752_wire_constant when (BITSEL_u32_u1_746_wire(0) /=  '0') else CONCAT_u4_u8_758_wire_constant;
    -- flow-through select operator MUX_773_inst
    wval_774 <= CONCAT_u32_u64_768_wire when (BITSEL_u32_u1_764_wire(0) /=  '0') else CONCAT_u32_u64_772_wire;
    -- flow-through slice operator slice_736_inst
    slice_736_wire <= write_pointer_buffer(31 downto 1);
    -- interlock type_cast_740_inst
    process(CONCAT_u31_u34_739_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 33 downto 0) := CONCAT_u31_u34_739_wire(33 downto 0);
      type_cast_740_wire <= tmp_var; -- 
    end process;
    -- binary operator ADD_u36_u36_731_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, type_cast_730_wire_constant, tmp_var);
      buffer_address_732 <= tmp_var; --
    end process;
    -- binary operator ADD_u36_u36_741_inst
    process(buffer_address_732, type_cast_740_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buffer_address_732, type_cast_740_wire, tmp_var);
      element_pair_address_742 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_746_inst
    process(write_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(write_pointer_buffer, konst_745_wire_constant, tmp_var);
      BITSEL_u32_u1_746_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_764_inst
    process(write_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(write_pointer_buffer, konst_763_wire_constant, tmp_var);
      BITSEL_u32_u1_764_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u31_u34_739_inst
    process(slice_736_wire) -- 
      variable tmp_var : std_logic_vector(33 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_736_wire, type_cast_738_wire_constant, tmp_var);
      CONCAT_u31_u34_739_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_768_inst
    process(type_cast_766_wire_constant, q_w_data_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_766_wire_constant, q_w_data_buffer, tmp_var);
      CONCAT_u32_u64_768_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_772_inst
    process(q_w_data_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(q_w_data_buffer, type_cast_771_wire_constant, tmp_var);
      CONCAT_u32_u64_772_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_788_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_788_call_req_0;
      call_stmt_788_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_788_call_req_1;
      call_stmt_788_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_781_wire_constant & type_cast_783_wire_constant & bmask_760 & element_pair_address_742 & wval_774;
      ignore_788 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end setQueueElement_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity setQueuePointers is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    wp : in  std_logic_vector(31 downto 0);
    rp : in  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity setQueuePointers;
architecture setQueuePointers_arch of setQueuePointers is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 100)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal wp_buffer :  std_logic_vector(31 downto 0);
  signal wp_update_enable: Boolean;
  signal rp_buffer :  std_logic_vector(31 downto 0);
  signal rp_update_enable: Boolean;
  -- output port buffer signals
  signal setQueuePointers_CP_564_start: Boolean;
  signal setQueuePointers_CP_564_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_464_call_ack_0 : boolean;
  signal call_stmt_464_call_req_0 : boolean;
  signal call_stmt_464_call_req_1 : boolean;
  signal call_stmt_464_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "setQueuePointers_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 100) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= wp;
  wp_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(99 downto 68) <= rp;
  rp_buffer <= in_buffer_data_out(99 downto 68);
  in_buffer_data_in(tag_length + 99 downto 100) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 99 downto 100);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  setQueuePointers_CP_564_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "setQueuePointers_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueuePointers_CP_564_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= setQueuePointers_CP_564_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueuePointers_CP_564_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  setQueuePointers_CP_564: Block -- control-path 
    signal setQueuePointers_CP_564_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    setQueuePointers_CP_564_elements(0) <= setQueuePointers_CP_564_start;
    setQueuePointers_CP_564_symbol <= setQueuePointers_CP_564_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_464/call_stmt_464_update_start_
      -- CP-element group 0: 	 call_stmt_464/call_stmt_464_sample_start_
      -- CP-element group 0: 	 call_stmt_464/call_stmt_464_Update/$entry
      -- CP-element group 0: 	 call_stmt_464/call_stmt_464_Sample/crr
      -- CP-element group 0: 	 call_stmt_464/call_stmt_464_Update/ccr
      -- CP-element group 0: 	 call_stmt_464/$entry
      -- CP-element group 0: 	 call_stmt_464/call_stmt_464_Sample/$entry
      -- CP-element group 0: 	 $entry
      -- 
    crr_577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_564_elements(0), ack => call_stmt_464_call_req_0); -- 
    ccr_582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_564_elements(0), ack => call_stmt_464_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_464/call_stmt_464_sample_completed_
      -- CP-element group 1: 	 call_stmt_464/call_stmt_464_Sample/cra
      -- CP-element group 1: 	 call_stmt_464/call_stmt_464_Sample/$exit
      -- 
    cra_578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_464_call_ack_0, ack => setQueuePointers_CP_564_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 call_stmt_464/call_stmt_464_update_completed_
      -- CP-element group 2: 	 call_stmt_464/call_stmt_464_Update/$exit
      -- CP-element group 2: 	 call_stmt_464/$exit
      -- CP-element group 2: 	 call_stmt_464/call_stmt_464_Update/cca
      -- CP-element group 2: 	 $exit
      -- 
    cca_583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_464_call_ack_1, ack => setQueuePointers_CP_564_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_459_wire : std_logic_vector(35 downto 0);
    signal CONCAT_u32_u64_462_wire : std_logic_vector(63 downto 0);
    signal NOT_u8_u8_456_wire_constant : std_logic_vector(7 downto 0);
    signal ignore_464 : std_logic_vector(63 downto 0);
    signal konst_458_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_451_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_453_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_456_wire_constant <= "11111111";
    konst_458_wire_constant <= "000000000000000000000000000000001000";
    type_cast_451_wire_constant <= "0";
    type_cast_453_wire_constant <= "0";
    -- binary operator ADD_u36_u36_459_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_458_wire_constant, tmp_var);
      ADD_u36_u36_459_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_462_inst
    process(wp_buffer, rp_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(wp_buffer, rp_buffer, tmp_var);
      CONCAT_u32_u64_462_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_464_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_464_call_req_0;
      call_stmt_464_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_464_call_req_1;
      call_stmt_464_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_451_wire_constant & type_cast_453_wire_constant & NOT_u8_u8_456_wire_constant & ADD_u36_u36_459_wire & CONCAT_u32_u64_462_wire;
      ignore_464 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end setQueuePointers_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity transmitEngineDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    FREE_Q : in std_logic_vector(35 downto 0);
    LAST_READ_TX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
    CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(1 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(1 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(11 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_reqs : out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_acks : in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_data : out  std_logic_vector(5 downto 0);
    getTxPacketPointerFromServer_call_tag  :  out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_reqs : out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_acks : in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_data : in   std_logic_vector(32 downto 0);
    getTxPacketPointerFromServer_return_tag :  in   std_logic_vector(0 downto 0);
    transmitPacket_call_reqs : out  std_logic_vector(0 downto 0);
    transmitPacket_call_acks : in   std_logic_vector(0 downto 0);
    transmitPacket_call_data : out  std_logic_vector(31 downto 0);
    transmitPacket_call_tag  :  out  std_logic_vector(0 downto 0);
    transmitPacket_return_reqs : out  std_logic_vector(0 downto 0);
    transmitPacket_return_acks : in   std_logic_vector(0 downto 0);
    transmitPacket_return_data : in   std_logic_vector(0 downto 0);
    transmitPacket_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity transmitEngineDaemon;
architecture transmitEngineDaemon_arch of transmitEngineDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal transmitEngineDaemon_CP_3075_start: Boolean;
  signal transmitEngineDaemon_CP_3075_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getTxPacketPointerFromServer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_index : in  std_logic_vector(5 downto 0);
      pkt_pointer : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(36 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(32 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component transmitPacket is -- 
    generic (tag_length : integer); 
    port ( -- 
      packet_pointer : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(145 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_call_acks : in   std_logic_vector(1 downto 0);
      accessMemory_call_data : out  std_logic_vector(219 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(3 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_return_acks : in   std_logic_vector(1 downto 0);
      accessMemory_return_data : in   std_logic_vector(127 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal ncount_1639_1569_buf_req_0 : boolean;
  signal ncount_1639_1569_buf_ack_0 : boolean;
  signal NOT_u1_u1_1590_inst_ack_1 : boolean;
  signal NOT_u1_u1_1590_inst_req_1 : boolean;
  signal W_pkt_pointer_1575_delayed_4_0_1600_inst_req_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_inst_ack_1 : boolean;
  signal W_pkt_pointer_1575_delayed_4_0_1600_inst_ack_1 : boolean;
  signal call_stmt_1609_call_ack_1 : boolean;
  signal phi_stmt_1565_req_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_inst_ack_1 : boolean;
  signal if_stmt_1545_branch_req_0 : boolean;
  signal phi_stmt_1565_req_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_inst_req_1 : boolean;
  signal ADD_u32_u32_1629_inst_ack_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_inst_req_0 : boolean;
  signal phi_stmt_1565_ack_0 : boolean;
  signal W_count_1596_delayed_14_0_1631_inst_ack_0 : boolean;
  signal if_stmt_1545_branch_ack_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_inst_ack_0 : boolean;
  signal call_stmt_1625_call_req_1 : boolean;
  signal if_stmt_1545_branch_ack_0 : boolean;
  signal call_stmt_1580_call_req_0 : boolean;
  signal call_stmt_1576_call_req_0 : boolean;
  signal ncount_1639_1569_buf_req_1 : boolean;
  signal W_count_1596_delayed_14_0_1631_inst_req_0 : boolean;
  signal call_stmt_1576_call_ack_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_inst_req_1 : boolean;
  signal call_stmt_1580_call_ack_0 : boolean;
  signal call_stmt_1609_call_req_1 : boolean;
  signal do_while_stmt_1553_branch_req_0 : boolean;
  signal NOT_u1_u1_1590_inst_ack_0 : boolean;
  signal NOT_u1_u1_1590_inst_req_0 : boolean;
  signal AND_u6_u6_1564_inst_ack_1 : boolean;
  signal ADD_u32_u32_1629_inst_req_1 : boolean;
  signal AND_u6_u6_1564_inst_req_1 : boolean;
  signal W_count_1588_delayed_14_0_1613_inst_ack_1 : boolean;
  signal call_stmt_1576_call_ack_1 : boolean;
  signal W_pkt_pointer_1575_delayed_4_0_1600_inst_ack_0 : boolean;
  signal W_pkt_pointer_1575_delayed_4_0_1600_inst_req_0 : boolean;
  signal W_count_1588_delayed_14_0_1613_inst_req_1 : boolean;
  signal call_stmt_1576_call_req_1 : boolean;
  signal call_stmt_1580_call_ack_1 : boolean;
  signal AND_u6_u6_1564_inst_ack_0 : boolean;
  signal call_stmt_1609_call_ack_0 : boolean;
  signal call_stmt_1609_call_req_0 : boolean;
  signal call_stmt_1580_call_req_1 : boolean;
  signal W_count_1588_delayed_14_0_1613_inst_ack_0 : boolean;
  signal AND_u6_u6_1564_inst_req_0 : boolean;
  signal W_count_1588_delayed_14_0_1613_inst_req_0 : boolean;
  signal call_stmt_1625_call_ack_0 : boolean;
  signal call_stmt_1625_call_req_0 : boolean;
  signal ncount_1639_1569_buf_ack_1 : boolean;
  signal W_count_1596_delayed_14_0_1631_inst_req_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_inst_ack_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_inst_req_0 : boolean;
  signal do_while_stmt_1553_branch_ack_0 : boolean;
  signal do_while_stmt_1553_branch_ack_1 : boolean;
  signal call_stmt_1625_call_ack_1 : boolean;
  signal ADD_u32_u32_1629_inst_ack_0 : boolean;
  signal ADD_u32_u32_1629_inst_req_0 : boolean;
  signal W_count_1596_delayed_14_0_1631_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "transmitEngineDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  transmitEngineDaemon_CP_3075_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "transmitEngineDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_3075_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_3075_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_3075_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  transmitEngineDaemon_CP_3075: Block -- control-path 
    signal transmitEngineDaemon_CP_3075_elements: BooleanArray(86 downto 0);
    -- 
  begin -- 
    transmitEngineDaemon_CP_3075_elements(0) <= transmitEngineDaemon_CP_3075_start;
    transmitEngineDaemon_CP_3075_symbol <= transmitEngineDaemon_CP_3075_elements(3);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 assign_stmt_1542/WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1542/WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_Sample/req
      -- CP-element group 0: 	 assign_stmt_1542/$entry
      -- CP-element group 0: 	 assign_stmt_1542/WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_sample_start_
      -- CP-element group 0: 	 $entry
      -- 
    req_3088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(0), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_1542/WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1542/WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_Sample/ack
      -- CP-element group 1: 	 assign_stmt_1542/WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_Update/$entry
      -- CP-element group 1: 	 assign_stmt_1542/WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1542/WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_Update/req
      -- CP-element group 1: 	 assign_stmt_1542/WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_update_start_
      -- 
    ack_3089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_inst_ack_0, ack => transmitEngineDaemon_CP_3075_elements(1)); -- 
    req_3093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(1), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_inst_req_1); -- 
    -- CP-element group 2:  branch  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	86 
    -- CP-element group 2:  members (10) 
      -- CP-element group 2: 	 assign_stmt_1542/WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_update_completed_
      -- CP-element group 2: 	 assign_stmt_1542/WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_Update/ack
      -- CP-element group 2: 	 assign_stmt_1542/$exit
      -- CP-element group 2: 	 assign_stmt_1542/WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1543/merge_stmt_1544__entry__
      -- CP-element group 2: 	 branch_block_stmt_1543/merge_stmt_1544__entry___PhiReq/$exit
      -- CP-element group 2: 	 branch_block_stmt_1543/merge_stmt_1544__entry___PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_1543/merge_stmt_1544_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_1543/branch_block_stmt_1543__entry__
      -- CP-element group 2: 	 branch_block_stmt_1543/$entry
      -- 
    ack_3094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_inst_ack_1, ack => transmitEngineDaemon_CP_3075_elements(2)); -- 
    -- CP-element group 3:  transition  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 $exit
      -- CP-element group 3: 	 branch_block_stmt_1543/$exit
      -- CP-element group 3: 	 branch_block_stmt_1543/branch_block_stmt_1543__exit__
      -- 
    transmitEngineDaemon_CP_3075_elements(3) <= false; 
    -- CP-element group 4:  transition  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	85 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	86 
    -- CP-element group 4:  members (4) 
      -- CP-element group 4: 	 branch_block_stmt_1543/do_while_stmt_1553__exit__
      -- CP-element group 4: 	 branch_block_stmt_1543/disable_loopback
      -- CP-element group 4: 	 branch_block_stmt_1543/disable_loopback_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_1543/disable_loopback_PhiReq/$exit
      -- 
    transmitEngineDaemon_CP_3075_elements(4) <= transmitEngineDaemon_CP_3075_elements(85);
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	86 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	86 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1543/if_stmt_1545_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_1543/if_stmt_1545_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_1543/not_enabled_yet_loopback
      -- CP-element group 5: 	 branch_block_stmt_1543/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_1543/not_enabled_yet_loopback_PhiReq/$exit
      -- 
    if_choice_transition_3167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1545_branch_ack_1, ack => transmitEngineDaemon_CP_3075_elements(5)); -- 
    -- CP-element group 6:  merge  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	86 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (4) 
      -- CP-element group 6: 	 branch_block_stmt_1543/do_while_stmt_1553__entry__
      -- CP-element group 6: 	 branch_block_stmt_1543/if_stmt_1545__exit__
      -- CP-element group 6: 	 branch_block_stmt_1543/if_stmt_1545_else_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_1543/if_stmt_1545_else_link/else_choice_transition
      -- 
    else_choice_transition_3171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1545_branch_ack_0, ack => transmitEngineDaemon_CP_3075_elements(6)); -- 
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_1543/do_while_stmt_1553/$entry
      -- CP-element group 7: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553__entry__
      -- 
    transmitEngineDaemon_CP_3075_elements(7) <= transmitEngineDaemon_CP_3075_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	85 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553__exit__
      -- 
    -- Element group transmitEngineDaemon_CP_3075_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1543/do_while_stmt_1553/loop_back
      -- 
    -- Element group transmitEngineDaemon_CP_3075_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	83 
    -- CP-element group 10: 	84 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1543/do_while_stmt_1553/condition_done
      -- CP-element group 10: 	 branch_block_stmt_1543/do_while_stmt_1553/loop_taken/$entry
      -- CP-element group 10: 	 branch_block_stmt_1543/do_while_stmt_1553/loop_exit/$entry
      -- 
    transmitEngineDaemon_CP_3075_elements(10) <= transmitEngineDaemon_CP_3075_elements(15);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	82 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1543/do_while_stmt_1553/loop_body_done
      -- 
    transmitEngineDaemon_CP_3075_elements(11) <= transmitEngineDaemon_CP_3075_elements(82);
    -- CP-element group 12:  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	29 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/back_edge_to_loop_body
      -- 
    transmitEngineDaemon_CP_3075_elements(12) <= transmitEngineDaemon_CP_3075_elements(9);
    -- CP-element group 13:  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	31 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/first_time_through_loop_body
      -- 
    transmitEngineDaemon_CP_3075_elements(13) <= transmitEngineDaemon_CP_3075_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	25 
    -- CP-element group 14: 	26 
    -- CP-element group 14: 	81 
    -- CP-element group 14: 	16 
    -- CP-element group 14: 	20 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1555_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/$entry
      -- CP-element group 14: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/loop_body_start
      -- 
    -- Element group transmitEngineDaemon_CP_3075_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	81 
    -- CP-element group 15: 	19 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/condition_evaluated
      -- 
    condition_evaluated_3187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(15), ack => do_while_stmt_1553_branch_req_0); -- 
    transmitEngineDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(81) & transmitEngineDaemon_CP_3075_elements(19);
      gj_transmitEngineDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	25 
    -- CP-element group 16: 	14 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	19 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	21 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/aggregated_phi_sample_req
      -- CP-element group 16: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1565_sample_start__ps
      -- 
    transmitEngineDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(25) & transmitEngineDaemon_CP_3075_elements(14) & transmitEngineDaemon_CP_3075_elements(19);
      gj_transmitEngineDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	27 
    -- CP-element group 17: 	23 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	47 
    -- CP-element group 17: 	51 
    -- CP-element group 17: 	71 
    -- CP-element group 17: 	75 
    -- CP-element group 17: 	82 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	25 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/aggregated_phi_sample_ack
      -- CP-element group 17: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1555_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1565_sample_completed_
      -- 
    transmitEngineDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(27) & transmitEngineDaemon_CP_3075_elements(23);
      gj_transmitEngineDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	26 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	22 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1565_update_start__ps
      -- CP-element group 18: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/aggregated_phi_update_req
      -- 
    transmitEngineDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(26) & transmitEngineDaemon_CP_3075_elements(20);
      gj_transmitEngineDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	24 
    -- CP-element group 19: 	28 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	16 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/aggregated_phi_update_ack
      -- 
    transmitEngineDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(24) & transmitEngineDaemon_CP_3075_elements(28);
      gj_transmitEngineDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	44 
    -- CP-element group 20: 	79 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1555_update_start_
      -- 
    transmitEngineDaemon_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(14) & transmitEngineDaemon_CP_3075_elements(44) & transmitEngineDaemon_CP_3075_elements(79);
      gj_transmitEngineDaemon_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/AND_u6_u6_1564_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/AND_u6_u6_1564_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/AND_u6_u6_1564_sample_start_
      -- 
    rr_3204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(21), ack => AND_u6_u6_1564_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(16) & transmitEngineDaemon_CP_3075_elements(23);
      gj_transmitEngineDaemon_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	18 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/AND_u6_u6_1564_Update/cr
      -- CP-element group 22: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/AND_u6_u6_1564_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/AND_u6_u6_1564_update_start_
      -- 
    cr_3209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(22), ack => AND_u6_u6_1564_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(18) & transmitEngineDaemon_CP_3075_elements(24);
      gj_transmitEngineDaemon_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	17 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	21 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/AND_u6_u6_1564_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/AND_u6_u6_1564_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/AND_u6_u6_1564_sample_completed_
      -- 
    ra_3205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_1564_inst_ack_0, ack => transmitEngineDaemon_CP_3075_elements(23)); -- 
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	42 
    -- CP-element group 24: 	78 
    -- CP-element group 24: 	19 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	22 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1555_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/AND_u6_u6_1564_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/AND_u6_u6_1564_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/AND_u6_u6_1564_update_completed_
      -- 
    ca_3210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_1564_inst_ack_1, ack => transmitEngineDaemon_CP_3075_elements(24)); -- 
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	14 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	49 
    -- CP-element group 25: 	53 
    -- CP-element group 25: 	73 
    -- CP-element group 25: 	77 
    -- CP-element group 25: 	17 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	16 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1565_sample_start_
      -- 
    transmitEngineDaemon_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(14) & transmitEngineDaemon_CP_3075_elements(49) & transmitEngineDaemon_CP_3075_elements(53) & transmitEngineDaemon_CP_3075_elements(73) & transmitEngineDaemon_CP_3075_elements(77) & transmitEngineDaemon_CP_3075_elements(17);
      gj_transmitEngineDaemon_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	14 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	64 
    -- CP-element group 26: 	72 
    -- CP-element group 26: 	76 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	18 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1565_update_start_
      -- 
    transmitEngineDaemon_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(14) & transmitEngineDaemon_CP_3075_elements(64) & transmitEngineDaemon_CP_3075_elements(72) & transmitEngineDaemon_CP_3075_elements(76);
      gj_transmitEngineDaemon_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	17 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1565_sample_completed__ps
      -- 
    -- Element group transmitEngineDaemon_CP_3075_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	70 
    -- CP-element group 28: 	74 
    -- CP-element group 28: 	62 
    -- CP-element group 28: 	19 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1565_update_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1565_update_completed_
      -- 
    -- Element group transmitEngineDaemon_CP_3075_elements(28) is bound as output of CP function.
    -- CP-element group 29:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	12 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1565_loopback_trigger
      -- 
    transmitEngineDaemon_CP_3075_elements(29) <= transmitEngineDaemon_CP_3075_elements(12);
    -- CP-element group 30:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1565_loopback_sample_req
      -- CP-element group 30: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1565_loopback_sample_req_ps
      -- 
    phi_stmt_1565_loopback_sample_req_3220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1565_loopback_sample_req_3220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(30), ack => phi_stmt_1565_req_1); -- 
    -- Element group transmitEngineDaemon_CP_3075_elements(30) is bound as output of CP function.
    -- CP-element group 31:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	13 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1565_entry_trigger
      -- 
    transmitEngineDaemon_CP_3075_elements(31) <= transmitEngineDaemon_CP_3075_elements(13);
    -- CP-element group 32:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1565_entry_sample_req
      -- CP-element group 32: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1565_entry_sample_req_ps
      -- 
    phi_stmt_1565_entry_sample_req_3223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1565_entry_sample_req_3223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(32), ack => phi_stmt_1565_req_0); -- 
    -- Element group transmitEngineDaemon_CP_3075_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1565_phi_mux_ack
      -- CP-element group 33: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/phi_stmt_1565_phi_mux_ack_ps
      -- 
    phi_stmt_1565_phi_mux_ack_3226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1565_ack_0, ack => transmitEngineDaemon_CP_3075_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/type_cast_1568_sample_start__ps
      -- CP-element group 34: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/type_cast_1568_sample_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/type_cast_1568_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/type_cast_1568_sample_start_
      -- 
    -- Element group transmitEngineDaemon_CP_3075_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (2) 
      -- CP-element group 35: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/type_cast_1568_update_start__ps
      -- CP-element group 35: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/type_cast_1568_update_start_
      -- 
    -- Element group transmitEngineDaemon_CP_3075_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/type_cast_1568_update_completed__ps
      -- 
    transmitEngineDaemon_CP_3075_elements(36) <= transmitEngineDaemon_CP_3075_elements(37);
    -- CP-element group 37:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	36 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/type_cast_1568_update_completed_
      -- 
    -- Element group transmitEngineDaemon_CP_3075_elements(37) is a control-delay.
    cp_element_37_delay: control_delay_element  generic map(name => " 37_delay", delay_value => 1)  port map(req => transmitEngineDaemon_CP_3075_elements(35), ack => transmitEngineDaemon_CP_3075_elements(37), clk => clk, reset =>reset);
    -- CP-element group 38:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/R_ncount_1569_Sample/req
      -- CP-element group 38: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/R_ncount_1569_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/R_ncount_1569_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/R_ncount_1569_sample_start__ps
      -- 
    req_3247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(38), ack => ncount_1639_1569_buf_req_0); -- 
    -- Element group transmitEngineDaemon_CP_3075_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/R_ncount_1569_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/R_ncount_1569_Update/req
      -- CP-element group 39: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/R_ncount_1569_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/R_ncount_1569_update_start__ps
      -- 
    req_3252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(39), ack => ncount_1639_1569_buf_req_1); -- 
    -- Element group transmitEngineDaemon_CP_3075_elements(39) is bound as output of CP function.
    -- CP-element group 40:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/R_ncount_1569_Sample/ack
      -- CP-element group 40: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/R_ncount_1569_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/R_ncount_1569_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/R_ncount_1569_sample_completed__ps
      -- 
    ack_3248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_1639_1569_buf_ack_0, ack => transmitEngineDaemon_CP_3075_elements(40)); -- 
    -- CP-element group 41:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (4) 
      -- CP-element group 41: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/R_ncount_1569_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/R_ncount_1569_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/R_ncount_1569_update_completed__ps
      -- CP-element group 41: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/R_ncount_1569_Update/ack
      -- 
    ack_3253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_1639_1569_buf_ack_1, ack => transmitEngineDaemon_CP_3075_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	24 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: 	69 
    -- CP-element group 42: 	61 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1576_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1576_Sample/crr
      -- CP-element group 42: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1576_sample_start_
      -- 
    crr_3262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(42), ack => call_stmt_1576_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(24) & transmitEngineDaemon_CP_3075_elements(44) & transmitEngineDaemon_CP_3075_elements(69) & transmitEngineDaemon_CP_3075_elements(61);
      gj_transmitEngineDaemon_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	48 
    -- CP-element group 43: 	52 
    -- CP-element group 43: 	69 
    -- CP-element group 43: 	56 
    -- CP-element group 43: 	61 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1576_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1576_Update/ccr
      -- CP-element group 43: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1576_update_start_
      -- 
    ccr_3267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(43), ack => call_stmt_1576_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(48) & transmitEngineDaemon_CP_3075_elements(52) & transmitEngineDaemon_CP_3075_elements(69) & transmitEngineDaemon_CP_3075_elements(56) & transmitEngineDaemon_CP_3075_elements(61);
      gj_transmitEngineDaemon_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: 	20 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1576_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1576_Sample/cra
      -- CP-element group 44: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1576_sample_completed_
      -- 
    cra_3263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1576_call_ack_0, ack => transmitEngineDaemon_CP_3075_elements(44)); -- 
    -- CP-element group 45:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: 	50 
    -- CP-element group 45: 	66 
    -- CP-element group 45: 	54 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1576_Update/cca
      -- CP-element group 45: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1576_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1576_update_completed_
      -- 
    cca_3268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1576_call_ack_1, ack => transmitEngineDaemon_CP_3075_elements(45)); -- 
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	48 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1580_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1580_Sample/crr
      -- CP-element group 46: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1580_sample_start_
      -- 
    crr_3276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(46), ack => call_stmt_1580_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(45) & transmitEngineDaemon_CP_3075_elements(48);
      gj_transmitEngineDaemon_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	17 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	68 
    -- CP-element group 47: 	60 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1580_update_start_
      -- CP-element group 47: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1580_Update/ccr
      -- CP-element group 47: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1580_Update/$entry
      -- 
    ccr_3281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(47), ack => call_stmt_1580_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(17) & transmitEngineDaemon_CP_3075_elements(68) & transmitEngineDaemon_CP_3075_elements(60);
      gj_transmitEngineDaemon_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	43 
    -- CP-element group 48: 	46 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1580_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1580_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1580_Sample/cra
      -- 
    cra_3277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1580_call_ack_0, ack => transmitEngineDaemon_CP_3075_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	66 
    -- CP-element group 49: 	58 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	25 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1580_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1580_Update/cca
      -- CP-element group 49: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1580_Update/$exit
      -- 
    cca_3282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1580_call_ack_1, ack => transmitEngineDaemon_CP_3075_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	45 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	52 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/NOT_u1_u1_1590_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/NOT_u1_u1_1590_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/NOT_u1_u1_1590_sample_start_
      -- 
    rr_3290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(50), ack => NOT_u1_u1_1590_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(45) & transmitEngineDaemon_CP_3075_elements(52);
      gj_transmitEngineDaemon_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	17 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	68 
    -- CP-element group 51: 	60 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/NOT_u1_u1_1590_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/NOT_u1_u1_1590_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/NOT_u1_u1_1590_update_start_
      -- 
    cr_3295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(51), ack => NOT_u1_u1_1590_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(17) & transmitEngineDaemon_CP_3075_elements(68) & transmitEngineDaemon_CP_3075_elements(60);
      gj_transmitEngineDaemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	43 
    -- CP-element group 52: 	50 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/NOT_u1_u1_1590_Sample/ra
      -- CP-element group 52: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/NOT_u1_u1_1590_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/NOT_u1_u1_1590_sample_completed_
      -- 
    ra_3291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1590_inst_ack_0, ack => transmitEngineDaemon_CP_3075_elements(52)); -- 
    -- CP-element group 53:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	66 
    -- CP-element group 53: 	58 
    -- CP-element group 53: marked-successors 
    -- CP-element group 53: 	25 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/NOT_u1_u1_1590_Update/ca
      -- CP-element group 53: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/NOT_u1_u1_1590_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/NOT_u1_u1_1590_update_completed_
      -- 
    ca_3296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1590_inst_ack_1, ack => transmitEngineDaemon_CP_3075_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	45 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1602_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1602_Sample/req
      -- CP-element group 54: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1602_Sample/$entry
      -- 
    req_3304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(54), ack => W_pkt_pointer_1575_delayed_4_0_1600_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(45) & transmitEngineDaemon_CP_3075_elements(56);
      gj_transmitEngineDaemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	60 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1602_Update/req
      -- CP-element group 55: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1602_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1602_update_start_
      -- 
    req_3309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(55), ack => W_pkt_pointer_1575_delayed_4_0_1600_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_3075_elements(60);
      gj_transmitEngineDaemon_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	43 
    -- CP-element group 56: 	54 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1602_Sample/ack
      -- CP-element group 56: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1602_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1602_sample_completed_
      -- 
    ack_3305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_pointer_1575_delayed_4_0_1600_inst_ack_0, ack => transmitEngineDaemon_CP_3075_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1602_Update/ack
      -- CP-element group 57: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1602_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1602_update_completed_
      -- 
    ack_3310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_pointer_1575_delayed_4_0_1600_inst_ack_1, ack => transmitEngineDaemon_CP_3075_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	49 
    -- CP-element group 58: 	53 
    -- CP-element group 58: 	57 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1609_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1609_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1609_Sample/crr
      -- 
    crr_3318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(58), ack => call_stmt_1609_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(49) & transmitEngineDaemon_CP_3075_elements(53) & transmitEngineDaemon_CP_3075_elements(57) & transmitEngineDaemon_CP_3075_elements(60);
      gj_transmitEngineDaemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1609_update_start_
      -- CP-element group 59: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1609_Update/ccr
      -- CP-element group 59: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1609_Update/$entry
      -- 
    ccr_3323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(59), ack => call_stmt_1609_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_3075_elements(61);
      gj_transmitEngineDaemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	47 
    -- CP-element group 60: 	51 
    -- CP-element group 60: 	55 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1609_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1609_Sample/cra
      -- CP-element group 60: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1609_Sample/$exit
      -- 
    cra_3319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1609_call_ack_0, ack => transmitEngineDaemon_CP_3075_elements(60)); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	82 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	42 
    -- CP-element group 61: 	43 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1609_Update/cca
      -- CP-element group 61: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1609_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1609_Update/$exit
      -- 
    cca_3324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1609_call_ack_1, ack => transmitEngineDaemon_CP_3075_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	28 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1615_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1615_Sample/req
      -- CP-element group 62: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1615_Sample/$entry
      -- 
    req_3332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(62), ack => W_count_1588_delayed_14_0_1613_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(28) & transmitEngineDaemon_CP_3075_elements(64);
      gj_transmitEngineDaemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	68 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1615_update_start_
      -- CP-element group 63: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1615_Update/req
      -- CP-element group 63: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1615_Update/$entry
      -- 
    req_3337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(63), ack => W_count_1588_delayed_14_0_1613_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_3075_elements(68);
      gj_transmitEngineDaemon_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	26 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1615_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1615_Sample/ack
      -- CP-element group 64: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1615_Sample/$exit
      -- 
    ack_3333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_1588_delayed_14_0_1613_inst_ack_0, ack => transmitEngineDaemon_CP_3075_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1615_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1615_Update/ack
      -- CP-element group 65: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1615_Update/$exit
      -- 
    ack_3338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_1588_delayed_14_0_1613_inst_ack_1, ack => transmitEngineDaemon_CP_3075_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	45 
    -- CP-element group 66: 	49 
    -- CP-element group 66: 	53 
    -- CP-element group 66: 	65 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1625_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1625_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1625_Sample/crr
      -- 
    crr_3346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(66), ack => call_stmt_1625_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(45) & transmitEngineDaemon_CP_3075_elements(49) & transmitEngineDaemon_CP_3075_elements(53) & transmitEngineDaemon_CP_3075_elements(65) & transmitEngineDaemon_CP_3075_elements(68);
      gj_transmitEngineDaemon_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1625_Update/ccr
      -- CP-element group 67: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1625_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1625_update_start_
      -- 
    ccr_3351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(67), ack => call_stmt_1625_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_3075_elements(69);
      gj_transmitEngineDaemon_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	47 
    -- CP-element group 68: 	51 
    -- CP-element group 68: 	63 
    -- CP-element group 68: 	66 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1625_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1625_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1625_Sample/cra
      -- 
    cra_3347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1625_call_ack_0, ack => transmitEngineDaemon_CP_3075_elements(68)); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	82 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	42 
    -- CP-element group 69: 	43 
    -- CP-element group 69: 	67 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1625_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1625_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/call_stmt_1625_Update/cca
      -- 
    cca_3352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1625_call_ack_1, ack => transmitEngineDaemon_CP_3075_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	28 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/ADD_u32_u32_1629_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/ADD_u32_u32_1629_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/ADD_u32_u32_1629_Sample/rr
      -- 
    rr_3360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(70), ack => ADD_u32_u32_1629_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(28) & transmitEngineDaemon_CP_3075_elements(72);
      gj_transmitEngineDaemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	17 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/ADD_u32_u32_1629_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/ADD_u32_u32_1629_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/ADD_u32_u32_1629_Update/$entry
      -- 
    cr_3365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(71), ack => ADD_u32_u32_1629_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(17) & transmitEngineDaemon_CP_3075_elements(73);
      gj_transmitEngineDaemon_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	26 
    -- CP-element group 72: 	70 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/ADD_u32_u32_1629_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/ADD_u32_u32_1629_Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/ADD_u32_u32_1629_Sample/$exit
      -- 
    ra_3361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_1629_inst_ack_0, ack => transmitEngineDaemon_CP_3075_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	82 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	25 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/ADD_u32_u32_1629_Update/ca
      -- CP-element group 73: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/ADD_u32_u32_1629_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/ADD_u32_u32_1629_Update/$exit
      -- 
    ca_3366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_1629_inst_ack_1, ack => transmitEngineDaemon_CP_3075_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	28 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1633_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1633_Sample/req
      -- CP-element group 74: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1633_sample_start_
      -- 
    req_3374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(74), ack => W_count_1596_delayed_14_0_1631_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(28) & transmitEngineDaemon_CP_3075_elements(76);
      gj_transmitEngineDaemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	17 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1633_update_start_
      -- CP-element group 75: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1633_Update/req
      -- CP-element group 75: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1633_Update/$entry
      -- 
    req_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(75), ack => W_count_1596_delayed_14_0_1631_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(17) & transmitEngineDaemon_CP_3075_elements(77);
      gj_transmitEngineDaemon_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	26 
    -- CP-element group 76: 	74 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1633_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1633_Sample/ack
      -- CP-element group 76: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1633_sample_completed_
      -- 
    ack_3375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_1596_delayed_14_0_1631_inst_ack_0, ack => transmitEngineDaemon_CP_3075_elements(76)); -- 
    -- CP-element group 77:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	82 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	25 
    -- CP-element group 77: 	75 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1633_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1633_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/assign_stmt_1633_Update/ack
      -- 
    ack_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_1596_delayed_14_0_1631_inst_ack_1, ack => transmitEngineDaemon_CP_3075_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	24 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	80 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_Sample/req
      -- CP-element group 78: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_Sample/$entry
      -- 
    req_3388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(78), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(24) & transmitEngineDaemon_CP_3075_elements(80);
      gj_transmitEngineDaemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	20 
    -- CP-element group 79:  members (6) 
      -- CP-element group 79: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_Update/req
      -- CP-element group 79: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_update_start_
      -- CP-element group 79: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_Sample/ack
      -- CP-element group 79: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_Sample/$exit
      -- 
    ack_3389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_inst_ack_0, ack => transmitEngineDaemon_CP_3075_elements(79)); -- 
    req_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(79), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_inst_req_1); -- 
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	78 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_Update/ack
      -- CP-element group 80: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_Update/$exit
      -- 
    ack_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_inst_ack_1, ack => transmitEngineDaemon_CP_3075_elements(80)); -- 
    -- CP-element group 81:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	14 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	15 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group transmitEngineDaemon_CP_3075_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => transmitEngineDaemon_CP_3075_elements(14), ack => transmitEngineDaemon_CP_3075_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  join  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	69 
    -- CP-element group 82: 	73 
    -- CP-element group 82: 	77 
    -- CP-element group 82: 	61 
    -- CP-element group 82: 	80 
    -- CP-element group 82: 	17 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	11 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1543/do_while_stmt_1553/do_while_stmt_1553_loop_body/$exit
      -- 
    transmitEngineDaemon_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 31,1 => 31,2 => 31,3 => 31,4 => 31,5 => 31);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3075_elements(69) & transmitEngineDaemon_CP_3075_elements(73) & transmitEngineDaemon_CP_3075_elements(77) & transmitEngineDaemon_CP_3075_elements(61) & transmitEngineDaemon_CP_3075_elements(80) & transmitEngineDaemon_CP_3075_elements(17);
      gj_transmitEngineDaemon_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	10 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1543/do_while_stmt_1553/loop_exit/$exit
      -- CP-element group 83: 	 branch_block_stmt_1543/do_while_stmt_1553/loop_exit/ack
      -- 
    ack_3399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1553_branch_ack_0, ack => transmitEngineDaemon_CP_3075_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	10 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1543/do_while_stmt_1553/loop_taken/$exit
      -- CP-element group 84: 	 branch_block_stmt_1543/do_while_stmt_1553/loop_taken/ack
      -- 
    ack_3403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1553_branch_ack_1, ack => transmitEngineDaemon_CP_3075_elements(84)); -- 
    -- CP-element group 85:  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	8 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	4 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1543/do_while_stmt_1553/$exit
      -- 
    transmitEngineDaemon_CP_3075_elements(85) <= transmitEngineDaemon_CP_3075_elements(8);
    -- CP-element group 86:  merge  branch  transition  place  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	2 
    -- CP-element group 86: 	4 
    -- CP-element group 86: 	5 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	5 
    -- CP-element group 86: 	6 
    -- CP-element group 86:  members (49) 
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/$entry
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/$exit
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/BITSEL_u32_u1_1548_inputs/RPIPE_CONTROL_REGISTER_1546/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/BITSEL_u32_u1_1548_inputs/RPIPE_CONTROL_REGISTER_1546/Update/ack
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/$entry
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/$exit
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/SplitProtocol/Update/ca
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/branch_req
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_if_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/BITSEL_u32_u1_1548_inputs/$entry
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_else_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/BITSEL_u32_u1_1548_inputs/$exit
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/BITSEL_u32_u1_1548_inputs/RPIPE_CONTROL_REGISTER_1546/$entry
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/BITSEL_u32_u1_1548_inputs/RPIPE_CONTROL_REGISTER_1546/$exit
      -- CP-element group 86: 	 branch_block_stmt_1543/NOT_u1_u1_1549_place
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/BITSEL_u32_u1_1548_inputs/RPIPE_CONTROL_REGISTER_1546/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/$exit
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/BITSEL_u32_u1_1548_inputs/RPIPE_CONTROL_REGISTER_1546/Update/req
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545__entry__
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/SplitProtocol/Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/$entry
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/SplitProtocol/Update/ca
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/BITSEL_u32_u1_1548_inputs/RPIPE_CONTROL_REGISTER_1546/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_1543/merge_stmt_1544__exit__
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/SplitProtocol/Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_dead_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/BITSEL_u32_u1_1548_inputs/RPIPE_CONTROL_REGISTER_1546/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_1543/merge_stmt_1544_PhiAck/$exit
      -- CP-element group 86: 	 branch_block_stmt_1543/merge_stmt_1544_PhiAck/dummy
      -- CP-element group 86: 	 branch_block_stmt_1543/merge_stmt_1544_PhiReqMerge
      -- CP-element group 86: 	 branch_block_stmt_1543/merge_stmt_1544_PhiAck/$entry
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/BITSEL_u32_u1_1548_inputs/RPIPE_CONTROL_REGISTER_1546/Sample/ack
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/BITSEL_u32_u1_1548_inputs/RPIPE_CONTROL_REGISTER_1546/Sample/req
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_1543/if_stmt_1545_eval_test/NOT_u1_u1_1549/BITSEL_u32_u1_1548/SplitProtocol/$exit
      -- 
    branch_req_3162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3075_elements(86), ack => if_stmt_1545_branch_req_0); -- 
    transmitEngineDaemon_CP_3075_elements(86) <= OrReduce(transmitEngineDaemon_CP_3075_elements(2) & transmitEngineDaemon_CP_3075_elements(4) & transmitEngineDaemon_CP_3075_elements(5));
    transmitEngineDaemon_do_while_stmt_1553_terminator_3404: loop_terminator -- 
      generic map (name => " transmitEngineDaemon_do_while_stmt_1553_terminator_3404", max_iterations_in_flight =>31) 
      port map(loop_body_exit => transmitEngineDaemon_CP_3075_elements(11),loop_continue => transmitEngineDaemon_CP_3075_elements(84),loop_terminate => transmitEngineDaemon_CP_3075_elements(83),loop_back => transmitEngineDaemon_CP_3075_elements(9),loop_exit => transmitEngineDaemon_CP_3075_elements(8),clk => clk, reset => reset); -- 
    phi_stmt_1565_phi_seq_3254_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitEngineDaemon_CP_3075_elements(31);
      transmitEngineDaemon_CP_3075_elements(34)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitEngineDaemon_CP_3075_elements(34);
      transmitEngineDaemon_CP_3075_elements(35)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitEngineDaemon_CP_3075_elements(36);
      transmitEngineDaemon_CP_3075_elements(32) <= phi_mux_reqs(0);
      triggers(1)  <= transmitEngineDaemon_CP_3075_elements(29);
      transmitEngineDaemon_CP_3075_elements(38)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitEngineDaemon_CP_3075_elements(40);
      transmitEngineDaemon_CP_3075_elements(39)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitEngineDaemon_CP_3075_elements(41);
      transmitEngineDaemon_CP_3075_elements(30) <= phi_mux_reqs(1);
      phi_stmt_1565_phi_seq_3254 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1565_phi_seq_3254") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitEngineDaemon_CP_3075_elements(16), 
          phi_sample_ack => transmitEngineDaemon_CP_3075_elements(27), 
          phi_update_req => transmitEngineDaemon_CP_3075_elements(18), 
          phi_update_ack => transmitEngineDaemon_CP_3075_elements(28), 
          phi_mux_ack => transmitEngineDaemon_CP_3075_elements(33), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3188_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= transmitEngineDaemon_CP_3075_elements(12);
        preds(1)  <= transmitEngineDaemon_CP_3075_elements(13);
        entry_tmerge_3188 : transition_merge -- 
          generic map(name => " entry_tmerge_3188")
          port map (preds => preds, symbol_out => transmitEngineDaemon_CP_3075_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_1595_1595_delayed_14_0_1630 : std_logic_vector(31 downto 0);
    signal ADD_u6_u6_1559_wire : std_logic_vector(5 downto 0);
    signal AND_u6_u6_1564_wire : std_logic_vector(5 downto 0);
    signal BITSEL_u32_u1_1548_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_1648_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1549_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1564_1564_delayed_4_0_1591 : std_logic_vector(0 downto 0);
    signal NOT_u4_u4_1621_wire_constant : std_logic_vector(3 downto 0);
    signal RPIPE_CONTROL_REGISTER_1546_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CONTROL_REGISTER_1646_wire : std_logic_vector(31 downto 0);
    signal RPIPE_FREE_Q_1606_wire : std_logic_vector(35 downto 0);
    signal RPIPE_LAST_READ_TX_QUEUE_INDEX_1557_wire : std_logic_vector(5 downto 0);
    signal RPIPE_NUMBER_OF_SERVERS_1560_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_1562_wire : std_logic_vector(31 downto 0);
    signal count_1565 : std_logic_vector(31 downto 0);
    signal count_1588_delayed_14_0_1615 : std_logic_vector(31 downto 0);
    signal count_1596_delayed_14_0_1633 : std_logic_vector(31 downto 0);
    signal ignore_resp_1625 : std_logic_vector(31 downto 0);
    signal konst_1541_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1547_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1558_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1561_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1622_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1628_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1647_wire_constant : std_logic_vector(31 downto 0);
    signal ncount_1639 : std_logic_vector(31 downto 0);
    signal ncount_1639_1569_buffered : std_logic_vector(31 downto 0);
    signal pkt_pointer_1575_delayed_4_0_1602 : std_logic_vector(31 downto 0);
    signal pkt_pointer_1576 : std_logic_vector(31 downto 0);
    signal push_pointer_back_to_free_Q_1596 : std_logic_vector(0 downto 0);
    signal push_status_1609 : std_logic_vector(0 downto 0);
    signal transmitted_flag_1580 : std_logic_vector(0 downto 0);
    signal tx_flag_1576 : std_logic_vector(0 downto 0);
    signal tx_q_index_1555 : std_logic_vector(5 downto 0);
    signal type_cast_1563_wire : std_logic_vector(5 downto 0);
    signal type_cast_1568_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1605_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1618_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_1621_wire_constant <= "1111";
    konst_1541_wire_constant <= "000000";
    konst_1547_wire_constant <= "00000000000000000000000000000000";
    konst_1558_wire_constant <= "000001";
    konst_1561_wire_constant <= "00000000000000000000000000000001";
    konst_1622_wire_constant <= "010101";
    konst_1628_wire_constant <= "00000000000000000000000000000001";
    konst_1647_wire_constant <= "00000000000000000000000000000000";
    type_cast_1568_wire_constant <= "00000000000000000000000000000001";
    type_cast_1605_wire_constant <= "1";
    type_cast_1618_wire_constant <= "0";
    phi_stmt_1565: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1568_wire_constant & ncount_1639_1569_buffered;
      req <= phi_stmt_1565_req_0 & phi_stmt_1565_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1565",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1565_ack_0,
          idata => idata,
          odata => count_1565,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1565
    -- flow-through select operator MUX_1638_inst
    ncount_1639 <= ADD_u32_u32_1595_1595_delayed_14_0_1630 when (push_pointer_back_to_free_Q_1596(0) /=  '0') else count_1596_delayed_14_0_1633;
    W_count_1588_delayed_14_0_1613_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_count_1588_delayed_14_0_1613_inst_req_0;
      W_count_1588_delayed_14_0_1613_inst_ack_0<= wack(0);
      rreq(0) <= W_count_1588_delayed_14_0_1613_inst_req_1;
      W_count_1588_delayed_14_0_1613_inst_ack_1<= rack(0);
      W_count_1588_delayed_14_0_1613_inst : InterlockBuffer generic map ( -- 
        name => "W_count_1588_delayed_14_0_1613_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_1565,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => count_1588_delayed_14_0_1615,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_count_1596_delayed_14_0_1631_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_count_1596_delayed_14_0_1631_inst_req_0;
      W_count_1596_delayed_14_0_1631_inst_ack_0<= wack(0);
      rreq(0) <= W_count_1596_delayed_14_0_1631_inst_req_1;
      W_count_1596_delayed_14_0_1631_inst_ack_1<= rack(0);
      W_count_1596_delayed_14_0_1631_inst : InterlockBuffer generic map ( -- 
        name => "W_count_1596_delayed_14_0_1631_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_1565,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => count_1596_delayed_14_0_1633,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_pkt_pointer_1575_delayed_4_0_1600_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_pkt_pointer_1575_delayed_4_0_1600_inst_req_0;
      W_pkt_pointer_1575_delayed_4_0_1600_inst_ack_0<= wack(0);
      rreq(0) <= W_pkt_pointer_1575_delayed_4_0_1600_inst_req_1;
      W_pkt_pointer_1575_delayed_4_0_1600_inst_ack_1<= rack(0);
      W_pkt_pointer_1575_delayed_4_0_1600_inst : InterlockBuffer generic map ( -- 
        name => "W_pkt_pointer_1575_delayed_4_0_1600_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => pkt_pointer_1576,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pkt_pointer_1575_delayed_4_0_1602,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    ncount_1639_1569_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ncount_1639_1569_buf_req_0;
      ncount_1639_1569_buf_ack_0<= wack(0);
      rreq(0) <= ncount_1639_1569_buf_req_1;
      ncount_1639_1569_buf_ack_1<= rack(0);
      ncount_1639_1569_buf : InterlockBuffer generic map ( -- 
        name => "ncount_1639_1569_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ncount_1639,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ncount_1639_1569_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1555
    process(AND_u6_u6_1564_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := AND_u6_u6_1564_wire(5 downto 0);
      tx_q_index_1555 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1563_inst
    process(SUB_u32_u32_1562_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := SUB_u32_u32_1562_wire(5 downto 0);
      type_cast_1563_wire <= tmp_var; -- 
    end process;
    do_while_stmt_1553_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_1648_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1553_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1553_branch_req_0,
          ack0 => do_while_stmt_1553_branch_ack_0,
          ack1 => do_while_stmt_1553_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1545_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1549_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1545_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1545_branch_req_0,
          ack0 => if_stmt_1545_branch_ack_0,
          ack1 => if_stmt_1545_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u32_u32_1629_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= count_1565;
      ADD_u32_u32_1595_1595_delayed_14_0_1630 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_1629_inst_req_0;
      ADD_u32_u32_1629_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_1629_inst_req_1;
      ADD_u32_u32_1629_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator ADD_u6_u6_1559_inst
    process(RPIPE_LAST_READ_TX_QUEUE_INDEX_1557_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(RPIPE_LAST_READ_TX_QUEUE_INDEX_1557_wire, konst_1558_wire_constant, tmp_var);
      ADD_u6_u6_1559_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1595_inst
    process(NOT_u1_u1_1564_1564_delayed_4_0_1591, transmitted_flag_1580) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_1564_1564_delayed_4_0_1591, transmitted_flag_1580, tmp_var);
      push_pointer_back_to_free_Q_1596 <= tmp_var; --
    end process;
    -- shared split operator group (3) : AND_u6_u6_1564_inst 
    ApIntAnd_group_3: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u6_u6_1559_wire & type_cast_1563_wire;
      AND_u6_u6_1564_wire <= data_out(5 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u6_u6_1564_inst_req_0;
      AND_u6_u6_1564_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u6_u6_1564_inst_req_1;
      AND_u6_u6_1564_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 6, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- binary operator BITSEL_u32_u1_1548_inst
    process(RPIPE_CONTROL_REGISTER_1546_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1546_wire, konst_1547_wire_constant, tmp_var);
      BITSEL_u32_u1_1548_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1648_inst
    process(RPIPE_CONTROL_REGISTER_1646_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1646_wire, konst_1647_wire_constant, tmp_var);
      BITSEL_u32_u1_1648_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1549_inst
    process(BITSEL_u32_u1_1548_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_1548_wire, tmp_var);
      NOT_u1_u1_1549_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (7) : NOT_u1_u1_1590_inst 
    ApIntNot_group_7: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= tx_flag_1576;
      NOT_u1_u1_1564_1564_delayed_4_0_1591 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1590_inst_req_0;
      NOT_u1_u1_1590_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1590_inst_req_1;
      NOT_u1_u1_1590_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_7_gI: SplitGuardInterface generic map(name => "ApIntNot_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- binary operator SUB_u32_u32_1562_inst
    process(RPIPE_NUMBER_OF_SERVERS_1560_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(RPIPE_NUMBER_OF_SERVERS_1560_wire, konst_1561_wire_constant, tmp_var);
      SUB_u32_u32_1562_wire <= tmp_var; --
    end process;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1546_wire <= CONTROL_REGISTER;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1646_wire <= CONTROL_REGISTER;
    -- read from input-signal FREE_Q
    RPIPE_FREE_Q_1606_wire <= FREE_Q;
    -- read from input-signal LAST_READ_TX_QUEUE_INDEX
    RPIPE_LAST_READ_TX_QUEUE_INDEX_1557_wire <= LAST_READ_TX_QUEUE_INDEX;
    -- read from input-signal NUMBER_OF_SERVERS
    RPIPE_NUMBER_OF_SERVERS_1560_wire <= NUMBER_OF_SERVERS;
    -- shared outport operator group (0) : WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_inst_req_0;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_inst_req_1;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_1540_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_1541_wire_constant;
      LAST_READ_TX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_READ_TX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_READ_TX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_READ_TX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(1),
          oack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(1),
          odata => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(11 downto 6),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_inst_req_0;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_inst_req_1;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_1642_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= tx_q_index_1555;
      LAST_READ_TX_QUEUE_INDEX_write_1_gI: SplitGuardInterface generic map(name => "LAST_READ_TX_QUEUE_INDEX_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_READ_TX_QUEUE_INDEX_write_1: OutputPortRevised -- 
        generic map ( name => "LAST_READ_TX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(5 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_1576_call 
    getTxPacketPointerFromServer_call_group_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(32 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 10);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1576_call_req_0;
      call_stmt_1576_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1576_call_req_1;
      call_stmt_1576_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getTxPacketPointerFromServer_call_group_0_gI: SplitGuardInterface generic map(name => "getTxPacketPointerFromServer_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tx_q_index_1555;
      pkt_pointer_1576 <= data_out(32 downto 1);
      tx_flag_1576 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 6,
        owidth => 6,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getTxPacketPointerFromServer_call_reqs(0),
          ackR => getTxPacketPointerFromServer_call_acks(0),
          dataR => getTxPacketPointerFromServer_call_data(5 downto 0),
          tagR => getTxPacketPointerFromServer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 33,
          owidth => 33,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getTxPacketPointerFromServer_return_acks(0), -- cross-over
          ackL => getTxPacketPointerFromServer_return_reqs(0), -- cross-over
          dataL => getTxPacketPointerFromServer_return_data(32 downto 0),
          tagL => getTxPacketPointerFromServer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1580_call 
    transmitPacket_call_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1580_call_req_0;
      call_stmt_1580_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1580_call_req_1;
      call_stmt_1580_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not tx_flag_1576(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      transmitPacket_call_group_1_gI: SplitGuardInterface generic map(name => "transmitPacket_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= pkt_pointer_1576;
      transmitted_flag_1580 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => transmitPacket_call_reqs(0),
          ackR => transmitPacket_call_acks(0),
          dataR => transmitPacket_call_data(31 downto 0),
          tagR => transmitPacket_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => transmitPacket_return_acks(0), -- cross-over
          ackL => transmitPacket_return_reqs(0), -- cross-over
          dataL => transmitPacket_return_data(0 downto 0),
          tagL => transmitPacket_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1609_call 
    pushIntoQueue_call_group_2: Block -- 
      signal data_in: std_logic_vector(68 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1609_call_req_0;
      call_stmt_1609_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1609_call_req_1;
      call_stmt_1609_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= push_pointer_back_to_free_Q_1596(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_2_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1605_wire_constant & RPIPE_FREE_Q_1606_wire & pkt_pointer_1575_delayed_4_0_1602;
      push_status_1609 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 69,
        owidth => 69,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(68 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_1625_call 
    AccessRegister_call_group_3: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1625_call_req_0;
      call_stmt_1625_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1625_call_req_1;
      call_stmt_1625_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= push_pointer_back_to_free_Q_1596(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_3_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1618_wire_constant & NOT_u4_u4_1621_wire_constant & konst_1622_wire_constant & count_1588_delayed_14_0_1615;
      ignore_resp_1625 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end transmitEngineDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity transmitPacket is -- 
  generic (tag_length : integer); 
  port ( -- 
    packet_pointer : in  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(1 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(1 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(145 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(1 downto 0);
    accessMemory_call_acks : in   std_logic_vector(1 downto 0);
    accessMemory_call_data : out  std_logic_vector(219 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(3 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(1 downto 0);
    accessMemory_return_acks : in   std_logic_vector(1 downto 0);
    accessMemory_return_data : in   std_logic_vector(127 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity transmitPacket;
architecture transmitPacket_arch of transmitPacket is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal packet_pointer_buffer :  std_logic_vector(31 downto 0);
  signal packet_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal transmitPacket_CP_2807_start: Boolean;
  signal transmitPacket_CP_2807_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal ncount_down_1488_1455_buf_ack_0 : boolean;
  signal SUB_u8_u8_1458_inst_req_0 : boolean;
  signal ncount_down_1488_1455_buf_req_1 : boolean;
  signal ADD_u36_u36_1463_inst_ack_0 : boolean;
  signal do_while_stmt_1451_branch_req_0 : boolean;
  signal phi_stmt_1459_req_1 : boolean;
  signal call_stmt_1438_call_ack_1 : boolean;
  signal ncount_down_1488_1455_buf_req_0 : boolean;
  signal phi_stmt_1459_req_0 : boolean;
  signal call_stmt_1438_call_ack_0 : boolean;
  signal phi_stmt_1459_ack_0 : boolean;
  signal ncount_down_1488_1455_buf_ack_1 : boolean;
  signal SUB_u8_u8_1458_inst_ack_0 : boolean;
  signal ADD_u36_u36_1463_inst_req_0 : boolean;
  signal ADD_u36_u36_1463_inst_ack_1 : boolean;
  signal SUB_u8_u8_1458_inst_req_1 : boolean;
  signal SUB_u8_u8_1458_inst_ack_1 : boolean;
  signal call_stmt_1438_call_req_0 : boolean;
  signal phi_stmt_1453_req_0 : boolean;
  signal phi_stmt_1453_req_1 : boolean;
  signal ADD_u36_u36_1463_inst_req_1 : boolean;
  signal call_stmt_1438_call_req_1 : boolean;
  signal phi_stmt_1453_ack_0 : boolean;
  signal nmem_addr_1493_1464_buf_req_0 : boolean;
  signal nmem_addr_1493_1464_buf_ack_0 : boolean;
  signal nmem_addr_1493_1464_buf_req_1 : boolean;
  signal nmem_addr_1493_1464_buf_ack_1 : boolean;
  signal call_stmt_1475_call_req_0 : boolean;
  signal call_stmt_1475_call_ack_0 : boolean;
  signal call_stmt_1475_call_req_1 : boolean;
  signal call_stmt_1475_call_ack_1 : boolean;
  signal CONCAT_u65_u73_1482_inst_req_0 : boolean;
  signal CONCAT_u65_u73_1482_inst_ack_0 : boolean;
  signal CONCAT_u65_u73_1482_inst_req_1 : boolean;
  signal CONCAT_u65_u73_1482_inst_ack_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1476_inst_req_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1476_inst_ack_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1476_inst_req_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1476_inst_ack_1 : boolean;
  signal do_while_stmt_1451_branch_ack_0 : boolean;
  signal do_while_stmt_1451_branch_ack_1 : boolean;
  signal call_stmt_1518_call_req_0 : boolean;
  signal call_stmt_1518_call_ack_0 : boolean;
  signal call_stmt_1518_call_req_1 : boolean;
  signal call_stmt_1518_call_ack_1 : boolean;
  signal CONCAT_u65_u73_1527_inst_req_0 : boolean;
  signal CONCAT_u65_u73_1527_inst_ack_0 : boolean;
  signal CONCAT_u65_u73_1527_inst_req_1 : boolean;
  signal CONCAT_u65_u73_1527_inst_ack_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1521_inst_req_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1521_inst_ack_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1521_inst_req_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1521_inst_ack_1 : boolean;
  signal EQ_u8_u1_1535_inst_req_0 : boolean;
  signal EQ_u8_u1_1535_inst_ack_0 : boolean;
  signal EQ_u8_u1_1535_inst_req_1 : boolean;
  signal EQ_u8_u1_1535_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "transmitPacket_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= packet_pointer;
  packet_pointer_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  transmitPacket_CP_2807_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "transmitPacket_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= status_buffer;
  status <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitPacket_CP_2807_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= transmitPacket_CP_2807_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitPacket_CP_2807_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  transmitPacket_CP_2807: Block -- control-path 
    signal transmitPacket_CP_2807_elements: BooleanArray(81 downto 0);
    -- 
  begin -- 
    transmitPacket_CP_2807_elements(0) <= transmitPacket_CP_2807_start;
    transmitPacket_CP_2807_symbol <= transmitPacket_CP_2807_elements(81);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_1425_to_assign_stmt_1446/call_stmt_1438_update_start_
      -- CP-element group 0: 	 assign_stmt_1425_to_assign_stmt_1446/call_stmt_1438_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1425_to_assign_stmt_1446/call_stmt_1438_sample_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_1425_to_assign_stmt_1446/call_stmt_1438_Sample/crr
      -- CP-element group 0: 	 assign_stmt_1425_to_assign_stmt_1446/call_stmt_1438_Update/ccr
      -- CP-element group 0: 	 assign_stmt_1425_to_assign_stmt_1446/call_stmt_1438_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1425_to_assign_stmt_1446/$entry
      -- 
    ccr_2825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(0), ack => call_stmt_1438_call_req_1); -- 
    crr_2820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(0), ack => call_stmt_1438_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_1425_to_assign_stmt_1446/call_stmt_1438_Sample/cra
      -- CP-element group 1: 	 assign_stmt_1425_to_assign_stmt_1446/call_stmt_1438_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1425_to_assign_stmt_1446/call_stmt_1438_sample_completed_
      -- 
    cra_2821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1438_call_ack_0, ack => transmitPacket_CP_2807_elements(1)); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (7) 
      -- CP-element group 2: 	 assign_stmt_1425_to_assign_stmt_1446/call_stmt_1438_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_1450/$entry
      -- CP-element group 2: 	 branch_block_stmt_1450/branch_block_stmt_1450__entry__
      -- CP-element group 2: 	 assign_stmt_1425_to_assign_stmt_1446/call_stmt_1438_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1450/do_while_stmt_1451__entry__
      -- CP-element group 2: 	 assign_stmt_1425_to_assign_stmt_1446/call_stmt_1438_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1425_to_assign_stmt_1446/$exit
      -- 
    cca_2826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1438_call_ack_1, ack => transmitPacket_CP_2807_elements(2)); -- 
    -- CP-element group 3:  fork  transition  place  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	72 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	74 
    -- CP-element group 3: 	73 
    -- CP-element group 3: 	79 
    -- CP-element group 3: 	80 
    -- CP-element group 3: 	76 
    -- CP-element group 3:  members (18) 
      -- CP-element group 3: 	 branch_block_stmt_1450/do_while_stmt_1451__exit__
      -- CP-element group 3: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536__entry__
      -- CP-element group 3: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/$entry
      -- CP-element group 3: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/call_stmt_1518_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/call_stmt_1518_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/call_stmt_1518_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/call_stmt_1518_Sample/crr
      -- CP-element group 3: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/call_stmt_1518_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/call_stmt_1518_Update/ccr
      -- CP-element group 3: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/CONCAT_u65_u73_1527_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/CONCAT_u65_u73_1527_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/CONCAT_u65_u73_1527_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/EQ_u8_u1_1535_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/EQ_u8_u1_1535_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/EQ_u8_u1_1535_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/EQ_u8_u1_1535_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/EQ_u8_u1_1535_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/EQ_u8_u1_1535_Update/cr
      -- 
    crr_3026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(3), ack => call_stmt_1518_call_req_0); -- 
    ccr_3031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(3), ack => call_stmt_1518_call_req_1); -- 
    cr_3045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(3), ack => CONCAT_u65_u73_1527_inst_req_1); -- 
    rr_3068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(3), ack => EQ_u8_u1_1535_inst_req_0); -- 
    cr_3073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(3), ack => EQ_u8_u1_1535_inst_req_1); -- 
    transmitPacket_CP_2807_elements(3) <= transmitPacket_CP_2807_elements(72);
    -- CP-element group 4:  transition  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_1450/do_while_stmt_1451/$entry
      -- CP-element group 4: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451__entry__
      -- 
    transmitPacket_CP_2807_elements(4) <= transmitPacket_CP_2807_elements(2);
    -- CP-element group 5:  merge  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	72 
    -- CP-element group 5:  members (1) 
      -- CP-element group 5: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451__exit__
      -- 
    -- Element group transmitPacket_CP_2807_elements(5) is bound as output of CP function.
    -- CP-element group 6:  merge  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1450/do_while_stmt_1451/loop_back
      -- 
    -- Element group transmitPacket_CP_2807_elements(6) is bound as output of CP function.
    -- CP-element group 7:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	70 
    -- CP-element group 7: 	71 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1450/do_while_stmt_1451/condition_done
      -- CP-element group 7: 	 branch_block_stmt_1450/do_while_stmt_1451/loop_exit/$entry
      -- CP-element group 7: 	 branch_block_stmt_1450/do_while_stmt_1451/loop_taken/$entry
      -- 
    transmitPacket_CP_2807_elements(7) <= transmitPacket_CP_2807_elements(12);
    -- CP-element group 8:  branch  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	69 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1450/do_while_stmt_1451/loop_body_done
      -- 
    transmitPacket_CP_2807_elements(8) <= transmitPacket_CP_2807_elements(69);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	23 
    -- CP-element group 9: 	42 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/back_edge_to_loop_body
      -- 
    transmitPacket_CP_2807_elements(9) <= transmitPacket_CP_2807_elements(6);
    -- CP-element group 10:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	44 
    -- CP-element group 10: 	25 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/first_time_through_loop_body
      -- 
    transmitPacket_CP_2807_elements(10) <= transmitPacket_CP_2807_elements(4);
    -- CP-element group 11:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	38 
    -- CP-element group 11: 	39 
    -- CP-element group 11: 	68 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	18 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/loop_body_start
      -- CP-element group 11: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/$entry
      -- 
    -- Element group transmitPacket_CP_2807_elements(11) is bound as output of CP function.
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	22 
    -- CP-element group 12: 	68 
    -- CP-element group 12: 	16 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	7 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/condition_evaluated
      -- 
    condition_evaluated_2850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(12), ack => do_while_stmt_1451_branch_req_0); -- 
    transmitPacket_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 31);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(22) & transmitPacket_CP_2807_elements(68) & transmitPacket_CP_2807_elements(16);
      gj_transmitPacket_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	17 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	19 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/aggregated_phi_sample_req
      -- CP-element group 13: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1459_sample_start__ps
      -- 
    transmitPacket_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(38) & transmitPacket_CP_2807_elements(17) & transmitPacket_CP_2807_elements(16);
      gj_transmitPacket_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	40 
    -- CP-element group 14: 	20 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	69 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	38 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1453_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1459_sample_completed_
      -- 
    transmitPacket_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(40) & transmitPacket_CP_2807_elements(20);
      gj_transmitPacket_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	39 
    -- CP-element group 15: 	18 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	21 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/aggregated_phi_update_req
      -- CP-element group 15: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1459_update_start__ps
      -- 
    transmitPacket_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(39) & transmitPacket_CP_2807_elements(18);
      gj_transmitPacket_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	41 
    -- CP-element group 16: 	22 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/aggregated_phi_update_ack
      -- 
    transmitPacket_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(41) & transmitPacket_CP_2807_elements(22);
      gj_transmitPacket_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	13 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1453_sample_start_
      -- 
    transmitPacket_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(11) & transmitPacket_CP_2807_elements(14);
      gj_transmitPacket_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	22 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	15 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1453_update_start_
      -- 
    transmitPacket_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(11) & transmitPacket_CP_2807_elements(22);
      gj_transmitPacket_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1453_sample_start__ps
      -- 
    transmitPacket_CP_2807_elements(19) <= transmitPacket_CP_2807_elements(13);
    -- CP-element group 20:  join  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1453_sample_completed__ps
      -- 
    -- Element group transmitPacket_CP_2807_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1453_update_start__ps
      -- 
    transmitPacket_CP_2807_elements(21) <= transmitPacket_CP_2807_elements(15);
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	12 
    -- CP-element group 22: 	16 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	18 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1453_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1453_update_completed__ps
      -- 
    -- Element group transmitPacket_CP_2807_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	9 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1453_loopback_trigger
      -- 
    transmitPacket_CP_2807_elements(23) <= transmitPacket_CP_2807_elements(9);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1453_loopback_sample_req
      -- CP-element group 24: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1453_loopback_sample_req_ps
      -- 
    phi_stmt_1453_loopback_sample_req_2865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1453_loopback_sample_req_2865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(24), ack => phi_stmt_1453_req_0); -- 
    -- Element group transmitPacket_CP_2807_elements(24) is bound as output of CP function.
    -- CP-element group 25:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	10 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1453_entry_trigger
      -- 
    transmitPacket_CP_2807_elements(25) <= transmitPacket_CP_2807_elements(10);
    -- CP-element group 26:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1453_entry_sample_req
      -- CP-element group 26: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1453_entry_sample_req_ps
      -- 
    phi_stmt_1453_entry_sample_req_2868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1453_entry_sample_req_2868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(26), ack => phi_stmt_1453_req_1); -- 
    -- Element group transmitPacket_CP_2807_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1453_phi_mux_ack
      -- CP-element group 27: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1453_phi_mux_ack_ps
      -- 
    phi_stmt_1453_phi_mux_ack_2871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1453_ack_0, ack => transmitPacket_CP_2807_elements(27)); -- 
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_ncount_down_1455_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_ncount_down_1455_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_ncount_down_1455_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_ncount_down_1455_sample_start_
      -- 
    req_2884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(28), ack => ncount_down_1488_1455_buf_req_0); -- 
    -- Element group transmitPacket_CP_2807_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_ncount_down_1455_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_ncount_down_1455_Update/req
      -- CP-element group 29: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_ncount_down_1455_update_start_
      -- CP-element group 29: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_ncount_down_1455_update_start__ps
      -- 
    req_2889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(29), ack => ncount_down_1488_1455_buf_req_1); -- 
    -- Element group transmitPacket_CP_2807_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_ncount_down_1455_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_ncount_down_1455_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_ncount_down_1455_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_ncount_down_1455_sample_completed__ps
      -- 
    ack_2885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_down_1488_1455_buf_ack_0, ack => transmitPacket_CP_2807_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_ncount_down_1455_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_ncount_down_1455_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_ncount_down_1455_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_ncount_down_1455_update_completed__ps
      -- 
    ack_2890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_down_1488_1455_buf_ack_1, ack => transmitPacket_CP_2807_elements(31)); -- 
    -- CP-element group 32:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/SUB_u8_u8_1458_sample_start__ps
      -- 
    -- Element group transmitPacket_CP_2807_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/SUB_u8_u8_1458_update_start__ps
      -- 
    -- Element group transmitPacket_CP_2807_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/SUB_u8_u8_1458_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/SUB_u8_u8_1458_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/SUB_u8_u8_1458_sample_start_
      -- 
    rr_2902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(34), ack => SUB_u8_u8_1458_inst_req_0); -- 
    transmitPacket_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(32) & transmitPacket_CP_2807_elements(36);
      gj_transmitPacket_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/SUB_u8_u8_1458_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/SUB_u8_u8_1458_Update/cr
      -- CP-element group 35: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/SUB_u8_u8_1458_update_start_
      -- 
    cr_2907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(35), ack => SUB_u8_u8_1458_inst_req_1); -- 
    transmitPacket_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(33) & transmitPacket_CP_2807_elements(37);
      gj_transmitPacket_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	34 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/SUB_u8_u8_1458_Sample/ra
      -- CP-element group 36: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/SUB_u8_u8_1458_sample_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/SUB_u8_u8_1458_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/SUB_u8_u8_1458_Sample/$exit
      -- 
    ra_2903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u8_u8_1458_inst_ack_0, ack => transmitPacket_CP_2807_elements(36)); -- 
    -- CP-element group 37:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	35 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/SUB_u8_u8_1458_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/SUB_u8_u8_1458_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/SUB_u8_u8_1458_Update/ca
      -- CP-element group 37: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/SUB_u8_u8_1458_update_completed__ps
      -- 
    ca_2908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u8_u8_1458_inst_ack_1, ack => transmitPacket_CP_2807_elements(37)); -- 
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	11 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	14 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	13 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1459_sample_start_
      -- 
    transmitPacket_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(11) & transmitPacket_CP_2807_elements(14);
      gj_transmitPacket_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	11 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	59 
    -- CP-element group 39: 	41 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	15 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1459_update_start_
      -- 
    transmitPacket_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(11) & transmitPacket_CP_2807_elements(59) & transmitPacket_CP_2807_elements(41);
      gj_transmitPacket_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	14 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1459_sample_completed__ps
      -- 
    -- Element group transmitPacket_CP_2807_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	57 
    -- CP-element group 41: 	16 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	39 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1459_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1459_update_completed__ps
      -- 
    -- Element group transmitPacket_CP_2807_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	9 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1459_loopback_trigger
      -- 
    transmitPacket_CP_2807_elements(42) <= transmitPacket_CP_2807_elements(9);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1459_loopback_sample_req_ps
      -- CP-element group 43: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1459_loopback_sample_req
      -- 
    phi_stmt_1459_loopback_sample_req_2919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1459_loopback_sample_req_2919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(43), ack => phi_stmt_1459_req_1); -- 
    -- Element group transmitPacket_CP_2807_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	10 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1459_entry_trigger
      -- 
    transmitPacket_CP_2807_elements(44) <= transmitPacket_CP_2807_elements(10);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1459_entry_sample_req_ps
      -- CP-element group 45: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1459_entry_sample_req
      -- 
    phi_stmt_1459_entry_sample_req_2922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1459_entry_sample_req_2922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(45), ack => phi_stmt_1459_req_0); -- 
    -- Element group transmitPacket_CP_2807_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1459_phi_mux_ack
      -- CP-element group 46: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/phi_stmt_1459_phi_mux_ack_ps
      -- 
    phi_stmt_1459_phi_mux_ack_2925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1459_ack_0, ack => transmitPacket_CP_2807_elements(46)); -- 
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/ADD_u36_u36_1463_sample_start__ps
      -- 
    -- Element group transmitPacket_CP_2807_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/ADD_u36_u36_1463_update_start__ps
      -- 
    -- Element group transmitPacket_CP_2807_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	51 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/ADD_u36_u36_1463_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/ADD_u36_u36_1463_Sample/rr
      -- CP-element group 49: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/ADD_u36_u36_1463_Sample/$entry
      -- 
    rr_2938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(49), ack => ADD_u36_u36_1463_inst_req_0); -- 
    transmitPacket_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(47) & transmitPacket_CP_2807_elements(51);
      gj_transmitPacket_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	52 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/ADD_u36_u36_1463_update_start_
      -- CP-element group 50: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/ADD_u36_u36_1463_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/ADD_u36_u36_1463_Update/cr
      -- 
    cr_2943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(50), ack => ADD_u36_u36_1463_inst_req_1); -- 
    transmitPacket_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(48) & transmitPacket_CP_2807_elements(52);
      gj_transmitPacket_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	49 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/ADD_u36_u36_1463_Sample/ra
      -- CP-element group 51: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/ADD_u36_u36_1463_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/ADD_u36_u36_1463_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/ADD_u36_u36_1463_sample_completed__ps
      -- 
    ra_2939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1463_inst_ack_0, ack => transmitPacket_CP_2807_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	50 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/ADD_u36_u36_1463_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/ADD_u36_u36_1463_update_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/ADD_u36_u36_1463_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/ADD_u36_u36_1463_update_completed_
      -- 
    ca_2944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1463_inst_ack_1, ack => transmitPacket_CP_2807_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_nmem_addr_1464_sample_start__ps
      -- CP-element group 53: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_nmem_addr_1464_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_nmem_addr_1464_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_nmem_addr_1464_Sample/req
      -- 
    req_2956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(53), ack => nmem_addr_1493_1464_buf_req_0); -- 
    -- Element group transmitPacket_CP_2807_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_nmem_addr_1464_update_start__ps
      -- CP-element group 54: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_nmem_addr_1464_update_start_
      -- CP-element group 54: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_nmem_addr_1464_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_nmem_addr_1464_Update/req
      -- 
    req_2961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(54), ack => nmem_addr_1493_1464_buf_req_1); -- 
    -- Element group transmitPacket_CP_2807_elements(54) is bound as output of CP function.
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_nmem_addr_1464_sample_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_nmem_addr_1464_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_nmem_addr_1464_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_nmem_addr_1464_Sample/ack
      -- 
    ack_2957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmem_addr_1493_1464_buf_ack_0, ack => transmitPacket_CP_2807_elements(55)); -- 
    -- CP-element group 56:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_nmem_addr_1464_update_completed__ps
      -- CP-element group 56: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_nmem_addr_1464_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_nmem_addr_1464_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/R_nmem_addr_1464_Update/ack
      -- 
    ack_2962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmem_addr_1493_1464_buf_ack_1, ack => transmitPacket_CP_2807_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	41 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	59 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/call_stmt_1475_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/call_stmt_1475_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/call_stmt_1475_Sample/crr
      -- 
    crr_2971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(57), ack => call_stmt_1475_call_req_0); -- 
    transmitPacket_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(41) & transmitPacket_CP_2807_elements(59);
      gj_transmitPacket_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	63 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/call_stmt_1475_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/call_stmt_1475_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/call_stmt_1475_Update/ccr
      -- 
    ccr_2976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(58), ack => call_stmt_1475_call_req_1); -- 
    transmitPacket_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(63) & transmitPacket_CP_2807_elements(60);
      gj_transmitPacket_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	39 
    -- CP-element group 59: 	57 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/call_stmt_1475_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/call_stmt_1475_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/call_stmt_1475_Sample/cra
      -- 
    cra_2972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1475_call_ack_0, ack => transmitPacket_CP_2807_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/call_stmt_1475_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/call_stmt_1475_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/call_stmt_1475_Update/cca
      -- 
    cca_2977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1475_call_ack_1, ack => transmitPacket_CP_2807_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/CONCAT_u65_u73_1482_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/CONCAT_u65_u73_1482_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/CONCAT_u65_u73_1482_Sample/rr
      -- 
    rr_2985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(61), ack => CONCAT_u65_u73_1482_inst_req_0); -- 
    transmitPacket_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(60) & transmitPacket_CP_2807_elements(63);
      gj_transmitPacket_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	66 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/CONCAT_u65_u73_1482_update_start_
      -- CP-element group 62: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/CONCAT_u65_u73_1482_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/CONCAT_u65_u73_1482_Update/cr
      -- 
    cr_2990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(62), ack => CONCAT_u65_u73_1482_inst_req_1); -- 
    transmitPacket_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(66) & transmitPacket_CP_2807_elements(64);
      gj_transmitPacket_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: 	58 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/CONCAT_u65_u73_1482_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/CONCAT_u65_u73_1482_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/CONCAT_u65_u73_1482_Sample/ra
      -- 
    ra_2986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_1482_inst_ack_0, ack => transmitPacket_CP_2807_elements(63)); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/CONCAT_u65_u73_1482_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/CONCAT_u65_u73_1482_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/CONCAT_u65_u73_1482_Update/ca
      -- 
    ca_2991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_1482_inst_ack_1, ack => transmitPacket_CP_2807_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/WPIPE_nic_to_mac_transmit_pipe_1476_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/WPIPE_nic_to_mac_transmit_pipe_1476_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/WPIPE_nic_to_mac_transmit_pipe_1476_Sample/req
      -- 
    req_2999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(65), ack => WPIPE_nic_to_mac_transmit_pipe_1476_inst_req_0); -- 
    transmitPacket_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(64) & transmitPacket_CP_2807_elements(67);
      gj_transmitPacket_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	62 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/WPIPE_nic_to_mac_transmit_pipe_1476_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/WPIPE_nic_to_mac_transmit_pipe_1476_update_start_
      -- CP-element group 66: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/WPIPE_nic_to_mac_transmit_pipe_1476_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/WPIPE_nic_to_mac_transmit_pipe_1476_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/WPIPE_nic_to_mac_transmit_pipe_1476_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/WPIPE_nic_to_mac_transmit_pipe_1476_Update/req
      -- 
    ack_3000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_1476_inst_ack_0, ack => transmitPacket_CP_2807_elements(66)); -- 
    req_3004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(66), ack => WPIPE_nic_to_mac_transmit_pipe_1476_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/WPIPE_nic_to_mac_transmit_pipe_1476_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/WPIPE_nic_to_mac_transmit_pipe_1476_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/WPIPE_nic_to_mac_transmit_pipe_1476_Update/ack
      -- 
    ack_3005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_1476_inst_ack_1, ack => transmitPacket_CP_2807_elements(67)); -- 
    -- CP-element group 68:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	11 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	12 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group transmitPacket_CP_2807_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => transmitPacket_CP_2807_elements(11), ack => transmitPacket_CP_2807_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	14 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	8 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1450/do_while_stmt_1451/do_while_stmt_1451_loop_body/$exit
      -- 
    transmitPacket_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(14) & transmitPacket_CP_2807_elements(67);
      gj_transmitPacket_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	7 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_1450/do_while_stmt_1451/loop_exit/$exit
      -- CP-element group 70: 	 branch_block_stmt_1450/do_while_stmt_1451/loop_exit/ack
      -- 
    ack_3010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1451_branch_ack_0, ack => transmitPacket_CP_2807_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	7 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_1450/do_while_stmt_1451/loop_taken/$exit
      -- CP-element group 71: 	 branch_block_stmt_1450/do_while_stmt_1451/loop_taken/ack
      -- 
    ack_3014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1451_branch_ack_1, ack => transmitPacket_CP_2807_elements(71)); -- 
    -- CP-element group 72:  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	5 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	3 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1450/do_while_stmt_1451/$exit
      -- 
    transmitPacket_CP_2807_elements(72) <= transmitPacket_CP_2807_elements(5);
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	3 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/call_stmt_1518_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/call_stmt_1518_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/call_stmt_1518_Sample/cra
      -- 
    cra_3027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1518_call_ack_0, ack => transmitPacket_CP_2807_elements(73)); -- 
    -- CP-element group 74:  transition  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	3 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (6) 
      -- CP-element group 74: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/call_stmt_1518_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/call_stmt_1518_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/call_stmt_1518_Update/cca
      -- CP-element group 74: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/CONCAT_u65_u73_1527_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/CONCAT_u65_u73_1527_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/CONCAT_u65_u73_1527_Sample/rr
      -- 
    cca_3032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1518_call_ack_1, ack => transmitPacket_CP_2807_elements(74)); -- 
    rr_3040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(74), ack => CONCAT_u65_u73_1527_inst_req_0); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/CONCAT_u65_u73_1527_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/CONCAT_u65_u73_1527_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/CONCAT_u65_u73_1527_Sample/ra
      -- 
    ra_3041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_1527_inst_ack_0, ack => transmitPacket_CP_2807_elements(75)); -- 
    -- CP-element group 76:  transition  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	3 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/CONCAT_u65_u73_1527_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/CONCAT_u65_u73_1527_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/CONCAT_u65_u73_1527_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/WPIPE_nic_to_mac_transmit_pipe_1521_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/WPIPE_nic_to_mac_transmit_pipe_1521_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/WPIPE_nic_to_mac_transmit_pipe_1521_Sample/req
      -- 
    ca_3046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_1527_inst_ack_1, ack => transmitPacket_CP_2807_elements(76)); -- 
    req_3054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(76), ack => WPIPE_nic_to_mac_transmit_pipe_1521_inst_req_0); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/WPIPE_nic_to_mac_transmit_pipe_1521_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/WPIPE_nic_to_mac_transmit_pipe_1521_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/WPIPE_nic_to_mac_transmit_pipe_1521_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/WPIPE_nic_to_mac_transmit_pipe_1521_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/WPIPE_nic_to_mac_transmit_pipe_1521_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/WPIPE_nic_to_mac_transmit_pipe_1521_Update/req
      -- 
    ack_3055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_1521_inst_ack_0, ack => transmitPacket_CP_2807_elements(77)); -- 
    req_3059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2807_elements(77), ack => WPIPE_nic_to_mac_transmit_pipe_1521_inst_req_1); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	81 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/WPIPE_nic_to_mac_transmit_pipe_1521_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/WPIPE_nic_to_mac_transmit_pipe_1521_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/WPIPE_nic_to_mac_transmit_pipe_1521_Update/ack
      -- 
    ack_3060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_1521_inst_ack_1, ack => transmitPacket_CP_2807_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	3 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/EQ_u8_u1_1535_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/EQ_u8_u1_1535_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/EQ_u8_u1_1535_Sample/ra
      -- 
    ra_3069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_1535_inst_ack_0, ack => transmitPacket_CP_2807_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	3 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/EQ_u8_u1_1535_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/EQ_u8_u1_1535_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/EQ_u8_u1_1535_Update/ca
      -- 
    ca_3074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_1535_inst_ack_1, ack => transmitPacket_CP_2807_elements(80)); -- 
    -- CP-element group 81:  join  transition  place  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: 	78 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536__exit__
      -- CP-element group 81: 	 branch_block_stmt_1450/$exit
      -- CP-element group 81: 	 $exit
      -- CP-element group 81: 	 branch_block_stmt_1450/branch_block_stmt_1450__exit__
      -- CP-element group 81: 	 branch_block_stmt_1450/call_stmt_1518_to_assign_stmt_1536/$exit
      -- 
    transmitPacket_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2807_elements(80) & transmitPacket_CP_2807_elements(78);
      gj_transmitPacket_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2807_elements(81), clk => clk, reset => reset); --
    end block;
    transmitPacket_do_while_stmt_1451_terminator_3015: loop_terminator -- 
      generic map (name => " transmitPacket_do_while_stmt_1451_terminator_3015", max_iterations_in_flight =>31) 
      port map(loop_body_exit => transmitPacket_CP_2807_elements(8),loop_continue => transmitPacket_CP_2807_elements(71),loop_terminate => transmitPacket_CP_2807_elements(70),loop_back => transmitPacket_CP_2807_elements(6),loop_exit => transmitPacket_CP_2807_elements(5),clk => clk, reset => reset); -- 
    phi_stmt_1453_phi_seq_2909_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitPacket_CP_2807_elements(23);
      transmitPacket_CP_2807_elements(28)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitPacket_CP_2807_elements(30);
      transmitPacket_CP_2807_elements(29)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitPacket_CP_2807_elements(31);
      transmitPacket_CP_2807_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= transmitPacket_CP_2807_elements(25);
      transmitPacket_CP_2807_elements(32)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitPacket_CP_2807_elements(36);
      transmitPacket_CP_2807_elements(33)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitPacket_CP_2807_elements(37);
      transmitPacket_CP_2807_elements(26) <= phi_mux_reqs(1);
      phi_stmt_1453_phi_seq_2909 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1453_phi_seq_2909") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitPacket_CP_2807_elements(19), 
          phi_sample_ack => transmitPacket_CP_2807_elements(20), 
          phi_update_req => transmitPacket_CP_2807_elements(21), 
          phi_update_ack => transmitPacket_CP_2807_elements(22), 
          phi_mux_ack => transmitPacket_CP_2807_elements(27), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1459_phi_seq_2963_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitPacket_CP_2807_elements(44);
      transmitPacket_CP_2807_elements(47)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitPacket_CP_2807_elements(51);
      transmitPacket_CP_2807_elements(48)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitPacket_CP_2807_elements(52);
      transmitPacket_CP_2807_elements(45) <= phi_mux_reqs(0);
      triggers(1)  <= transmitPacket_CP_2807_elements(42);
      transmitPacket_CP_2807_elements(53)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitPacket_CP_2807_elements(55);
      transmitPacket_CP_2807_elements(54)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitPacket_CP_2807_elements(56);
      transmitPacket_CP_2807_elements(43) <= phi_mux_reqs(1);
      phi_stmt_1459_phi_seq_2963 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1459_phi_seq_2963") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitPacket_CP_2807_elements(13), 
          phi_sample_ack => transmitPacket_CP_2807_elements(40), 
          phi_update_req => transmitPacket_CP_2807_elements(15), 
          phi_update_ack => transmitPacket_CP_2807_elements(41), 
          phi_mux_ack => transmitPacket_CP_2807_elements(46), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2851_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= transmitPacket_CP_2807_elements(9);
        preds(1)  <= transmitPacket_CP_2807_elements(10);
        entry_tmerge_2851 : transition_merge -- 
          generic map(name => " entry_tmerge_2851")
          port map (preds => preds, symbol_out => transmitPacket_CP_2807_elements(11));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_1463_wire : std_logic_vector(35 downto 0);
    signal CONCAT_u1_u65_1480_wire : std_logic_vector(64 downto 0);
    signal CONCAT_u1_u65_1525_wire : std_logic_vector(64 downto 0);
    signal CONCAT_u32_u36_1423_wire : std_logic_vector(35 downto 0);
    signal CONCAT_u65_u73_1482_wire : std_logic_vector(72 downto 0);
    signal CONCAT_u65_u73_1527_wire : std_logic_vector(72 downto 0);
    signal R_FULL_BYTE_MASK_1433_wire_constant : std_logic_vector(7 downto 0);
    signal R_FULL_BYTE_MASK_1470_wire_constant : std_logic_vector(7 downto 0);
    signal R_FULL_BYTE_MASK_1481_wire_constant : std_logic_vector(7 downto 0);
    signal R_FULL_BYTE_MASK_1513_wire_constant : std_logic_vector(7 downto 0);
    signal SUB_u36_u36_1533_wire : std_logic_vector(35 downto 0);
    signal SUB_u8_u8_1458_wire : std_logic_vector(7 downto 0);
    signal control_data_1438 : std_logic_vector(63 downto 0);
    signal control_data_addr_1425 : std_logic_vector(35 downto 0);
    signal count_down_1453 : std_logic_vector(7 downto 0);
    signal data_1475 : std_logic_vector(63 downto 0);
    signal konst_1457_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1462_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1486_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1491_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1502_wire_constant : std_logic_vector(7 downto 0);
    signal last_tkeep_1446 : std_logic_vector(7 downto 0);
    signal last_word_1518 : std_logic_vector(63 downto 0);
    signal mem_addr_1459 : std_logic_vector(35 downto 0);
    signal ncount_down_1488 : std_logic_vector(7 downto 0);
    signal ncount_down_1488_1455_buffered : std_logic_vector(7 downto 0);
    signal nmem_addr_1493 : std_logic_vector(35 downto 0);
    signal nmem_addr_1493_1464_buffered : std_logic_vector(35 downto 0);
    signal not_last_word_1504 : std_logic_vector(0 downto 0);
    signal packet_size_1442 : std_logic_vector(7 downto 0);
    signal slice_1420_wire : std_logic_vector(31 downto 0);
    signal type_cast_1422_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_1430_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1432_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1436_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1467_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1469_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1473_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1478_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1510_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1512_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1516_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1523_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1534_wire : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_FULL_BYTE_MASK_1433_wire_constant <= "11111111";
    R_FULL_BYTE_MASK_1470_wire_constant <= "11111111";
    R_FULL_BYTE_MASK_1481_wire_constant <= "11111111";
    R_FULL_BYTE_MASK_1513_wire_constant <= "11111111";
    konst_1457_wire_constant <= "00010000";
    konst_1462_wire_constant <= "000000000000000000000000000000011000";
    konst_1486_wire_constant <= "00001000";
    konst_1491_wire_constant <= "000000000000000000000000000000001000";
    konst_1502_wire_constant <= "00001000";
    type_cast_1422_wire_constant <= "0000";
    type_cast_1430_wire_constant <= "0";
    type_cast_1432_wire_constant <= "1";
    type_cast_1436_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1467_wire_constant <= "0";
    type_cast_1469_wire_constant <= "1";
    type_cast_1473_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1478_wire_constant <= "0";
    type_cast_1510_wire_constant <= "0";
    type_cast_1512_wire_constant <= "1";
    type_cast_1516_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1523_wire_constant <= "1";
    phi_stmt_1453: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ncount_down_1488_1455_buffered & SUB_u8_u8_1458_wire;
      req <= phi_stmt_1453_req_0 & phi_stmt_1453_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1453",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1453_ack_0,
          idata => idata,
          odata => count_down_1453,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1453
    phi_stmt_1459: Block -- phi operator 
      signal idata: std_logic_vector(71 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u36_u36_1463_wire & nmem_addr_1493_1464_buffered;
      req <= phi_stmt_1459_req_0 & phi_stmt_1459_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1459",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 36) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1459_ack_0,
          idata => idata,
          odata => mem_addr_1459,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1459
    -- flow-through slice operator slice_1420_inst
    slice_1420_wire <= packet_pointer_buffer(31 downto 0);
    -- flow-through slice operator slice_1441_inst
    packet_size_1442 <= control_data_1438(15 downto 8);
    -- flow-through slice operator slice_1445_inst
    last_tkeep_1446 <= control_data_1438(7 downto 0);
    ncount_down_1488_1455_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ncount_down_1488_1455_buf_req_0;
      ncount_down_1488_1455_buf_ack_0<= wack(0);
      rreq(0) <= ncount_down_1488_1455_buf_req_1;
      ncount_down_1488_1455_buf_ack_1<= rack(0);
      ncount_down_1488_1455_buf : InterlockBuffer generic map ( -- 
        name => "ncount_down_1488_1455_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ncount_down_1488,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ncount_down_1488_1455_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmem_addr_1493_1464_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmem_addr_1493_1464_buf_req_0;
      nmem_addr_1493_1464_buf_ack_0<= wack(0);
      rreq(0) <= nmem_addr_1493_1464_buf_req_1;
      nmem_addr_1493_1464_buf_ack_1<= rack(0);
      nmem_addr_1493_1464_buf : InterlockBuffer generic map ( -- 
        name => "nmem_addr_1493_1464_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmem_addr_1493,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmem_addr_1493_1464_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1424_inst
    process(CONCAT_u32_u36_1423_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 35 downto 0) := CONCAT_u32_u36_1423_wire(35 downto 0);
      control_data_addr_1425 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1534_inst
    process(SUB_u36_u36_1533_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := SUB_u36_u36_1533_wire(7 downto 0);
      type_cast_1534_wire <= tmp_var; -- 
    end process;
    do_while_stmt_1451_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= not_last_word_1504;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1451_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1451_branch_req_0,
          ack0 => do_while_stmt_1451_branch_ack_0,
          ack1 => do_while_stmt_1451_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u36_u36_1463_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= control_data_addr_1425;
      ADD_u36_u36_1463_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_1463_inst_req_0;
      ADD_u36_u36_1463_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_1463_inst_req_1;
      ADD_u36_u36_1463_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000011000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator ADD_u36_u36_1492_inst
    process(mem_addr_1459) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mem_addr_1459, konst_1491_wire_constant, tmp_var);
      nmem_addr_1493 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u65_1480_inst
    process(type_cast_1478_wire_constant, data_1475) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1478_wire_constant, data_1475, tmp_var);
      CONCAT_u1_u65_1480_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u65_1525_inst
    process(type_cast_1523_wire_constant, last_word_1518) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1523_wire_constant, last_word_1518, tmp_var);
      CONCAT_u1_u65_1525_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u36_1423_inst
    process(slice_1420_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1420_wire, type_cast_1422_wire_constant, tmp_var);
      CONCAT_u32_u36_1423_wire <= tmp_var; --
    end process;
    -- shared split operator group (5) : CONCAT_u65_u73_1482_inst 
    ApConcat_group_5: Block -- 
      signal data_in: std_logic_vector(64 downto 0);
      signal data_out: std_logic_vector(72 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u1_u65_1480_wire;
      CONCAT_u65_u73_1482_wire <= data_out(72 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u65_u73_1482_inst_req_0;
      CONCAT_u65_u73_1482_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u65_u73_1482_inst_req_1;
      CONCAT_u65_u73_1482_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_5_gI: SplitGuardInterface generic map(name => "ApConcat_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 65,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 73,
          constant_operand => "11111111",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : CONCAT_u65_u73_1527_inst 
    ApConcat_group_6: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal data_out: std_logic_vector(72 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u1_u65_1525_wire & last_tkeep_1446;
      CONCAT_u65_u73_1527_wire <= data_out(72 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u65_u73_1527_inst_req_0;
      CONCAT_u65_u73_1527_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u65_u73_1527_inst_req_1;
      CONCAT_u65_u73_1527_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_6_gI: SplitGuardInterface generic map(name => "ApConcat_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 65,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 73,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : EQ_u8_u1_1535_inst 
    ApIntEq_group_7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= packet_size_1442 & type_cast_1534_wire;
      status_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_1535_inst_req_0;
      EQ_u8_u1_1535_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_1535_inst_req_1;
      EQ_u8_u1_1535_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_7_gI: SplitGuardInterface generic map(name => "ApIntEq_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- binary operator SUB_u36_u36_1533_inst
    process(nmem_addr_1493, control_data_addr_1425) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntSub_proc(nmem_addr_1493, control_data_addr_1425, tmp_var);
      SUB_u36_u36_1533_wire <= tmp_var; --
    end process;
    -- shared split operator group (9) : SUB_u8_u8_1458_inst 
    ApIntSub_group_9: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= packet_size_1442;
      SUB_u8_u8_1458_wire <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u8_u8_1458_inst_req_0;
      SUB_u8_u8_1458_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u8_u8_1458_inst_req_1;
      SUB_u8_u8_1458_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_9_gI: SplitGuardInterface generic map(name => "ApIntSub_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00010000",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- binary operator SUB_u8_u8_1487_inst
    process(count_down_1453) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSub_proc(count_down_1453, konst_1486_wire_constant, tmp_var);
      ncount_down_1488 <= tmp_var; --
    end process;
    -- binary operator UGT_u8_u1_1503_inst
    process(ncount_down_1488) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ncount_down_1488, konst_1502_wire_constant, tmp_var);
      not_last_word_1504 <= tmp_var; --
    end process;
    -- shared outport operator group (0) : WPIPE_nic_to_mac_transmit_pipe_1476_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_1476_inst_req_0;
      WPIPE_nic_to_mac_transmit_pipe_1476_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_1476_inst_req_1;
      WPIPE_nic_to_mac_transmit_pipe_1476_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u65_u73_1482_wire;
      nic_to_mac_transmit_pipe_write_0_gI: SplitGuardInterface generic map(name => "nic_to_mac_transmit_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_to_mac_transmit_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "nic_to_mac_transmit_pipe", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_to_mac_transmit_pipe_pipe_write_req(1),
          oack => nic_to_mac_transmit_pipe_pipe_write_ack(1),
          odata => nic_to_mac_transmit_pipe_pipe_write_data(145 downto 73),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_nic_to_mac_transmit_pipe_1521_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_1521_inst_req_0;
      WPIPE_nic_to_mac_transmit_pipe_1521_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_1521_inst_req_1;
      WPIPE_nic_to_mac_transmit_pipe_1521_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u65_u73_1527_wire;
      nic_to_mac_transmit_pipe_write_1_gI: SplitGuardInterface generic map(name => "nic_to_mac_transmit_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_to_mac_transmit_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "nic_to_mac_transmit_pipe", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_to_mac_transmit_pipe_pipe_write_req(0),
          oack => nic_to_mac_transmit_pipe_pipe_write_ack(0),
          odata => nic_to_mac_transmit_pipe_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_1438_call call_stmt_1518_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(219 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1438_call_req_0;
      reqL_unguarded(0) <= call_stmt_1518_call_req_0;
      call_stmt_1438_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1518_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1438_call_req_1;
      reqR_unguarded(0) <= call_stmt_1518_call_req_1;
      call_stmt_1438_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1518_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1430_wire_constant & type_cast_1432_wire_constant & R_FULL_BYTE_MASK_1433_wire_constant & control_data_addr_1425 & type_cast_1436_wire_constant & type_cast_1510_wire_constant & type_cast_1512_wire_constant & R_FULL_BYTE_MASK_1513_wire_constant & nmem_addr_1493 & type_cast_1516_wire_constant;
      control_data_1438 <= data_out(127 downto 64);
      last_word_1518 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 220,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(1),
          ackR => accessMemory_call_acks(1),
          dataR => accessMemory_call_data(219 downto 110),
          tagR => accessMemory_call_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(1), -- cross-over
          ackL => accessMemory_return_reqs(1), -- cross-over
          dataL => accessMemory_return_data(127 downto 64),
          tagL => accessMemory_return_tag(3 downto 2),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1475_call 
    accessMemory_call_group_1: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 3);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1475_call_req_0;
      call_stmt_1475_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1475_call_req_1;
      call_stmt_1475_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_1_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1467_wire_constant & type_cast_1469_wire_constant & R_FULL_BYTE_MASK_1470_wire_constant & mem_addr_1459 & type_cast_1473_wire_constant;
      data_1475 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end transmitPacket_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity writeControlInformationToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    base_buffer_pointer : in  std_logic_vector(35 downto 0);
    packet_size : in  std_logic_vector(7 downto 0);
    last_keep : in  std_logic_vector(7 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeControlInformationToMem;
architecture writeControlInformationToMem_arch of writeControlInformationToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 52)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal base_buffer_pointer_buffer :  std_logic_vector(35 downto 0);
  signal base_buffer_pointer_update_enable: Boolean;
  signal packet_size_buffer :  std_logic_vector(7 downto 0);
  signal packet_size_update_enable: Boolean;
  signal last_keep_buffer :  std_logic_vector(7 downto 0);
  signal last_keep_update_enable: Boolean;
  -- output port buffer signals
  signal writeControlInformationToMem_CP_999_start: Boolean;
  signal writeControlInformationToMem_CP_999_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_694_call_ack_0 : boolean;
  signal call_stmt_694_call_ack_1 : boolean;
  signal call_stmt_694_call_req_1 : boolean;
  signal call_stmt_694_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeControlInformationToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 52) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= base_buffer_pointer;
  base_buffer_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(43 downto 36) <= packet_size;
  packet_size_buffer <= in_buffer_data_out(43 downto 36);
  in_buffer_data_in(51 downto 44) <= last_keep;
  last_keep_buffer <= in_buffer_data_out(51 downto 44);
  in_buffer_data_in(tag_length + 51 downto 52) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 51 downto 52);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeControlInformationToMem_CP_999_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeControlInformationToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_999_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_999_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_999_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeControlInformationToMem_CP_999: Block -- control-path 
    signal writeControlInformationToMem_CP_999_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    writeControlInformationToMem_CP_999_elements(0) <= writeControlInformationToMem_CP_999_start;
    writeControlInformationToMem_CP_999_symbol <= writeControlInformationToMem_CP_999_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_685_to_call_stmt_694/call_stmt_694_Update/$entry
      -- CP-element group 0: 	 assign_stmt_685_to_call_stmt_694/call_stmt_694_Update/ccr
      -- CP-element group 0: 	 assign_stmt_685_to_call_stmt_694/call_stmt_694_Sample/crr
      -- CP-element group 0: 	 assign_stmt_685_to_call_stmt_694/call_stmt_694_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_685_to_call_stmt_694/call_stmt_694_update_start_
      -- CP-element group 0: 	 assign_stmt_685_to_call_stmt_694/call_stmt_694_sample_start_
      -- CP-element group 0: 	 assign_stmt_685_to_call_stmt_694/$entry
      -- CP-element group 0: 	 $entry
      -- 
    crr_1012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeControlInformationToMem_CP_999_elements(0), ack => call_stmt_694_call_req_0); -- 
    ccr_1017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeControlInformationToMem_CP_999_elements(0), ack => call_stmt_694_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_685_to_call_stmt_694/call_stmt_694_Sample/cra
      -- CP-element group 1: 	 assign_stmt_685_to_call_stmt_694/call_stmt_694_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_685_to_call_stmt_694/call_stmt_694_sample_completed_
      -- 
    cra_1013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_694_call_ack_0, ack => writeControlInformationToMem_CP_999_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 assign_stmt_685_to_call_stmt_694/call_stmt_694_Update/$exit
      -- CP-element group 2: 	 assign_stmt_685_to_call_stmt_694/call_stmt_694_Update/cca
      -- CP-element group 2: 	 assign_stmt_685_to_call_stmt_694/call_stmt_694_update_completed_
      -- CP-element group 2: 	 assign_stmt_685_to_call_stmt_694/$exit
      -- CP-element group 2: 	 $exit
      -- 
    cca_1018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_694_call_ack_1, ack => writeControlInformationToMem_CP_999_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u8_u16_683_wire : std_logic_vector(15 downto 0);
    signal R_FULL_BYTE_MASK_690_wire_constant : std_logic_vector(7 downto 0);
    signal control_data_685 : std_logic_vector(63 downto 0);
    signal ignore_return_694 : std_logic_vector(63 downto 0);
    signal type_cast_687_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_689_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_FULL_BYTE_MASK_690_wire_constant <= "11111111";
    type_cast_687_wire_constant <= "0";
    type_cast_689_wire_constant <= "0";
    -- interlock type_cast_684_inst
    process(CONCAT_u8_u16_683_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := CONCAT_u8_u16_683_wire(15 downto 0);
      control_data_685 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_683_inst
    process(packet_size_buffer, last_keep_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(packet_size_buffer, last_keep_buffer, tmp_var);
      CONCAT_u8_u16_683_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_694_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_694_call_req_0;
      call_stmt_694_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_694_call_req_1;
      call_stmt_694_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_687_wire_constant & type_cast_689_wire_constant & R_FULL_BYTE_MASK_690_wire_constant & base_buffer_pointer_buffer & control_data_685;
      ignore_return_694 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writeControlInformationToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity writeEthernetHeaderToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    buf_pointer : in  std_logic_vector(35 downto 0);
    buf_position : out  std_logic_vector(35 downto 0);
    nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeEthernetHeaderToMem;
architecture writeEthernetHeaderToMem_arch of writeEthernetHeaderToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal buf_pointer_buffer :  std_logic_vector(35 downto 0);
  signal buf_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal buf_position_buffer :  std_logic_vector(35 downto 0);
  signal buf_position_update_enable: Boolean;
  signal writeEthernetHeaderToMem_CP_700_start: Boolean;
  signal writeEthernetHeaderToMem_CP_700_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal do_while_stmt_547_branch_req_0 : boolean;
  signal phi_stmt_549_req_1 : boolean;
  signal phi_stmt_549_req_0 : boolean;
  signal phi_stmt_549_ack_0 : boolean;
  signal ADD_u36_u36_553_inst_req_0 : boolean;
  signal ADD_u36_u36_553_inst_ack_0 : boolean;
  signal ADD_u36_u36_553_inst_req_1 : boolean;
  signal ADD_u36_u36_553_inst_ack_1 : boolean;
  signal nbuf_position_593_554_buf_req_0 : boolean;
  signal nbuf_position_593_554_buf_ack_0 : boolean;
  signal nbuf_position_593_554_buf_req_1 : boolean;
  signal nbuf_position_593_554_buf_ack_1 : boolean;
  signal phi_stmt_555_req_1 : boolean;
  signal phi_stmt_555_req_0 : boolean;
  signal phi_stmt_555_ack_0 : boolean;
  signal nI_588_559_buf_req_0 : boolean;
  signal nI_588_559_buf_ack_0 : boolean;
  signal nI_588_559_buf_req_1 : boolean;
  signal nI_588_559_buf_ack_1 : boolean;
  signal RPIPE_nic_rx_to_header_562_inst_req_0 : boolean;
  signal RPIPE_nic_rx_to_header_562_inst_ack_0 : boolean;
  signal RPIPE_nic_rx_to_header_562_inst_req_1 : boolean;
  signal RPIPE_nic_rx_to_header_562_inst_ack_1 : boolean;
  signal call_stmt_583_call_req_0 : boolean;
  signal call_stmt_583_call_ack_0 : boolean;
  signal call_stmt_583_call_req_1 : boolean;
  signal call_stmt_583_call_ack_1 : boolean;
  signal do_while_stmt_547_branch_ack_0 : boolean;
  signal do_while_stmt_547_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeEthernetHeaderToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= buf_pointer;
  buf_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeEthernetHeaderToMem_CP_700_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeEthernetHeaderToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 36) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(35 downto 0) <= buf_position_buffer;
  buf_position <= out_buffer_data_out(35 downto 0);
  out_buffer_data_in(tag_length + 35 downto 36) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 35 downto 36);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_700_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_700_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_700_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeEthernetHeaderToMem_CP_700: Block -- control-path 
    signal writeEthernetHeaderToMem_CP_700_elements: BooleanArray(66 downto 0);
    -- 
  begin -- 
    writeEthernetHeaderToMem_CP_700_elements(0) <= writeEthernetHeaderToMem_CP_700_start;
    writeEthernetHeaderToMem_CP_700_symbol <= writeEthernetHeaderToMem_CP_700_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_546/$entry
      -- CP-element group 0: 	 branch_block_stmt_546/branch_block_stmt_546__entry__
      -- CP-element group 0: 	 branch_block_stmt_546/do_while_stmt_547__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	66 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_546/$exit
      -- CP-element group 1: 	 branch_block_stmt_546/branch_block_stmt_546__exit__
      -- CP-element group 1: 	 branch_block_stmt_546/do_while_stmt_547__exit__
      -- 
    writeEthernetHeaderToMem_CP_700_elements(1) <= writeEthernetHeaderToMem_CP_700_elements(66);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_546/do_while_stmt_547/$entry
      -- CP-element group 2: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547__entry__
      -- 
    writeEthernetHeaderToMem_CP_700_elements(2) <= writeEthernetHeaderToMem_CP_700_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	66 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547__exit__
      -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_546/do_while_stmt_547/loop_back
      -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	64 
    -- CP-element group 5: 	65 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_546/do_while_stmt_547/condition_done
      -- CP-element group 5: 	 branch_block_stmt_546/do_while_stmt_547/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_546/do_while_stmt_547/loop_taken/$entry
      -- 
    writeEthernetHeaderToMem_CP_700_elements(5) <= writeEthernetHeaderToMem_CP_700_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	63 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_546/do_while_stmt_547/loop_body_done
      -- 
    writeEthernetHeaderToMem_CP_700_elements(6) <= writeEthernetHeaderToMem_CP_700_elements(63);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	40 
    -- CP-element group 7: 	21 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/back_edge_to_loop_body
      -- 
    writeEthernetHeaderToMem_CP_700_elements(7) <= writeEthernetHeaderToMem_CP_700_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	42 
    -- CP-element group 8: 	23 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/first_time_through_loop_body
      -- 
    writeEthernetHeaderToMem_CP_700_elements(8) <= writeEthernetHeaderToMem_CP_700_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	36 
    -- CP-element group 9: 	37 
    -- CP-element group 9: 	62 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	53 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_560_sample_start_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	62 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/condition_evaluated
      -- 
    condition_evaluated_724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_700_elements(10), ack => do_while_stmt_547_branch_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_700_elements(62) & writeEthernetHeaderToMem_CP_700_elements(14);
      gj_writeEthernetHeaderToMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_700_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	54 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_555_sample_start__ps
      -- 
    writeEthernetHeaderToMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_700_elements(36) & writeEthernetHeaderToMem_CP_700_elements(9) & writeEthernetHeaderToMem_CP_700_elements(15) & writeEthernetHeaderToMem_CP_700_elements(14);
      gj_writeEthernetHeaderToMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_700_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	38 
    -- CP-element group 12: 	56 
    -- CP-element group 12: 	18 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	63 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	36 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_549_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_555_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_560_sample_completed_
      -- 
    writeEthernetHeaderToMem_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_700_elements(38) & writeEthernetHeaderToMem_CP_700_elements(56) & writeEthernetHeaderToMem_CP_700_elements(18);
      gj_writeEthernetHeaderToMem_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_700_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	37 
    -- CP-element group 13: 	53 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	55 
    -- CP-element group 13: 	19 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_555_update_start__ps
      -- 
    writeEthernetHeaderToMem_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_700_elements(37) & writeEthernetHeaderToMem_CP_700_elements(53) & writeEthernetHeaderToMem_CP_700_elements(16);
      gj_writeEthernetHeaderToMem_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_700_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	57 
    -- CP-element group 14: 	20 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/aggregated_phi_update_ack
      -- 
    writeEthernetHeaderToMem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_700_elements(39) & writeEthernetHeaderToMem_CP_700_elements(57) & writeEthernetHeaderToMem_CP_700_elements(20);
      gj_writeEthernetHeaderToMem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_700_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_549_sample_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_700_elements(9) & writeEthernetHeaderToMem_CP_700_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_700_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_549_update_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_700_elements(9) & writeEthernetHeaderToMem_CP_700_elements(20);
      gj_writeEthernetHeaderToMem_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_700_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_549_sample_start__ps
      -- 
    writeEthernetHeaderToMem_CP_700_elements(17) <= writeEthernetHeaderToMem_CP_700_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_549_sample_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_549_update_start__ps
      -- 
    writeEthernetHeaderToMem_CP_700_elements(19) <= writeEthernetHeaderToMem_CP_700_elements(13);
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_549_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_549_update_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_549_loopback_trigger
      -- 
    writeEthernetHeaderToMem_CP_700_elements(21) <= writeEthernetHeaderToMem_CP_700_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_549_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_549_loopback_sample_req_ps
      -- 
    phi_stmt_549_loopback_sample_req_739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_549_loopback_sample_req_739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_700_elements(22), ack => phi_stmt_549_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_549_entry_trigger
      -- 
    writeEthernetHeaderToMem_CP_700_elements(23) <= writeEthernetHeaderToMem_CP_700_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_549_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_549_entry_sample_req_ps
      -- 
    phi_stmt_549_entry_sample_req_742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_549_entry_sample_req_742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_700_elements(24), ack => phi_stmt_549_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_549_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_549_phi_mux_ack_ps
      -- 
    phi_stmt_549_phi_mux_ack_745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_549_ack_0, ack => writeEthernetHeaderToMem_CP_700_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/ADD_u36_u36_553_sample_start__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/ADD_u36_u36_553_update_start__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/ADD_u36_u36_553_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/ADD_u36_u36_553_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/ADD_u36_u36_553_Sample/rr
      -- 
    rr_758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_700_elements(28), ack => ADD_u36_u36_553_inst_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_700_elements(26) & writeEthernetHeaderToMem_CP_700_elements(30);
      gj_writeEthernetHeaderToMem_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_700_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	31 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/ADD_u36_u36_553_update_start_
      -- CP-element group 29: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/ADD_u36_u36_553_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/ADD_u36_u36_553_Update/cr
      -- 
    cr_763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_700_elements(29), ack => ADD_u36_u36_553_inst_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_700_elements(27) & writeEthernetHeaderToMem_CP_700_elements(31);
      gj_writeEthernetHeaderToMem_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_700_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/ADD_u36_u36_553_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/ADD_u36_u36_553_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/ADD_u36_u36_553_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/ADD_u36_u36_553_Sample/ra
      -- 
    ra_759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_553_inst_ack_0, ack => writeEthernetHeaderToMem_CP_700_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: marked-successors 
    -- CP-element group 31: 	29 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/ADD_u36_u36_553_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/ADD_u36_u36_553_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/ADD_u36_u36_553_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/ADD_u36_u36_553_Update/ca
      -- 
    ca_764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_553_inst_ack_1, ack => writeEthernetHeaderToMem_CP_700_elements(31)); -- 
    -- CP-element group 32:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nbuf_position_554_sample_start__ps
      -- CP-element group 32: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nbuf_position_554_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nbuf_position_554_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nbuf_position_554_Sample/req
      -- 
    req_776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_700_elements(32), ack => nbuf_position_593_554_buf_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nbuf_position_554_update_start__ps
      -- CP-element group 33: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nbuf_position_554_update_start_
      -- CP-element group 33: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nbuf_position_554_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nbuf_position_554_Update/req
      -- 
    req_781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_700_elements(33), ack => nbuf_position_593_554_buf_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nbuf_position_554_sample_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nbuf_position_554_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nbuf_position_554_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nbuf_position_554_Sample/ack
      -- 
    ack_777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nbuf_position_593_554_buf_ack_0, ack => writeEthernetHeaderToMem_CP_700_elements(34)); -- 
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nbuf_position_554_update_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nbuf_position_554_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nbuf_position_554_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nbuf_position_554_Update/ack
      -- 
    ack_782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nbuf_position_593_554_buf_ack_1, ack => writeEthernetHeaderToMem_CP_700_elements(35)); -- 
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	9 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	12 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	11 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_555_sample_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_700_elements(9) & writeEthernetHeaderToMem_CP_700_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_700_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	9 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	13 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_555_update_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_700_elements(9) & writeEthernetHeaderToMem_CP_700_elements(39);
      gj_writeEthernetHeaderToMem_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_700_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	12 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_555_sample_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(38) is bound as output of CP function.
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_555_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_555_update_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_555_loopback_trigger
      -- 
    writeEthernetHeaderToMem_CP_700_elements(40) <= writeEthernetHeaderToMem_CP_700_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_555_loopback_sample_req
      -- CP-element group 41: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_555_loopback_sample_req_ps
      -- 
    phi_stmt_555_loopback_sample_req_793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_555_loopback_sample_req_793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_700_elements(41), ack => phi_stmt_555_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_555_entry_trigger
      -- 
    writeEthernetHeaderToMem_CP_700_elements(42) <= writeEthernetHeaderToMem_CP_700_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_555_entry_sample_req
      -- CP-element group 43: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_555_entry_sample_req_ps
      -- 
    phi_stmt_555_entry_sample_req_796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_555_entry_sample_req_796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_700_elements(43), ack => phi_stmt_555_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_555_phi_mux_ack
      -- CP-element group 44: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_555_phi_mux_ack_ps
      -- 
    phi_stmt_555_phi_mux_ack_799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_555_ack_0, ack => writeEthernetHeaderToMem_CP_700_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/type_cast_558_sample_start__ps
      -- CP-element group 45: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/type_cast_558_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/type_cast_558_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/type_cast_558_sample_completed_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/type_cast_558_update_start__ps
      -- CP-element group 46: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/type_cast_558_update_start_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/type_cast_558_update_completed__ps
      -- 
    writeEthernetHeaderToMem_CP_700_elements(47) <= writeEthernetHeaderToMem_CP_700_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/type_cast_558_update_completed_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => writeEthernetHeaderToMem_CP_700_elements(46), ack => writeEthernetHeaderToMem_CP_700_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nI_559_sample_start__ps
      -- CP-element group 49: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nI_559_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nI_559_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nI_559_Sample/req
      -- 
    req_820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_700_elements(49), ack => nI_588_559_buf_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nI_559_update_start__ps
      -- CP-element group 50: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nI_559_update_start_
      -- CP-element group 50: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nI_559_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nI_559_Update/req
      -- 
    req_825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_700_elements(50), ack => nI_588_559_buf_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nI_559_sample_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nI_559_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nI_559_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nI_559_Sample/ack
      -- 
    ack_821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_588_559_buf_ack_0, ack => writeEthernetHeaderToMem_CP_700_elements(51)); -- 
    -- CP-element group 52:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nI_559_update_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nI_559_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nI_559_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/R_nI_559_Update/ack
      -- 
    ack_826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_588_559_buf_ack_1, ack => writeEthernetHeaderToMem_CP_700_elements(52)); -- 
    -- CP-element group 53:  join  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	9 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	60 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	13 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_560_update_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_700_elements(9) & writeEthernetHeaderToMem_CP_700_elements(60);
      gj_writeEthernetHeaderToMem_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_700_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	11 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	57 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/RPIPE_nic_rx_to_header_562_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/RPIPE_nic_rx_to_header_562_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/RPIPE_nic_rx_to_header_562_Sample/rr
      -- 
    rr_839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_700_elements(54), ack => RPIPE_nic_rx_to_header_562_inst_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_700_elements(11) & writeEthernetHeaderToMem_CP_700_elements(57);
      gj_writeEthernetHeaderToMem_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_700_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	13 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/RPIPE_nic_rx_to_header_562_update_start_
      -- CP-element group 55: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/RPIPE_nic_rx_to_header_562_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/RPIPE_nic_rx_to_header_562_Update/cr
      -- 
    cr_844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_700_elements(55), ack => RPIPE_nic_rx_to_header_562_inst_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_700_elements(56) & writeEthernetHeaderToMem_CP_700_elements(13);
      gj_writeEthernetHeaderToMem_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_700_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: 	12 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/RPIPE_nic_rx_to_header_562_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/RPIPE_nic_rx_to_header_562_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/RPIPE_nic_rx_to_header_562_Sample/ra
      -- 
    ra_840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_header_562_inst_ack_0, ack => writeEthernetHeaderToMem_CP_700_elements(56)); -- 
    -- CP-element group 57:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	14 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	54 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/phi_stmt_560_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/RPIPE_nic_rx_to_header_562_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/RPIPE_nic_rx_to_header_562_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/RPIPE_nic_rx_to_header_562_Update/ca
      -- 
    ca_845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_header_562_inst_ack_1, ack => writeEthernetHeaderToMem_CP_700_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/call_stmt_583_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/call_stmt_583_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/call_stmt_583_Sample/crr
      -- 
    crr_853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_700_elements(58), ack => call_stmt_583_call_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_700_elements(57) & writeEthernetHeaderToMem_CP_700_elements(60);
      gj_writeEthernetHeaderToMem_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_700_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/call_stmt_583_update_start_
      -- CP-element group 59: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/call_stmt_583_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/call_stmt_583_Update/ccr
      -- 
    ccr_858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_700_elements(59), ack => call_stmt_583_call_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeEthernetHeaderToMem_CP_700_elements(61);
      gj_writeEthernetHeaderToMem_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_700_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: 	53 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/call_stmt_583_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/call_stmt_583_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/call_stmt_583_Sample/cra
      -- 
    cra_854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_583_call_ack_0, ack => writeEthernetHeaderToMem_CP_700_elements(60)); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/call_stmt_583_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/call_stmt_583_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/call_stmt_583_Update/cca
      -- 
    cca_859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_583_call_ack_1, ack => writeEthernetHeaderToMem_CP_700_elements(61)); -- 
    -- CP-element group 62:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	9 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	10 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group writeEthernetHeaderToMem_CP_700_elements(62) is a control-delay.
    cp_element_62_delay: control_delay_element  generic map(name => " 62_delay", delay_value => 1)  port map(req => writeEthernetHeaderToMem_CP_700_elements(9), ack => writeEthernetHeaderToMem_CP_700_elements(62), clk => clk, reset =>reset);
    -- CP-element group 63:  join  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: 	12 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	6 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_546/do_while_stmt_547/do_while_stmt_547_loop_body/$exit
      -- 
    writeEthernetHeaderToMem_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_700_elements(61) & writeEthernetHeaderToMem_CP_700_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_700_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	5 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_546/do_while_stmt_547/loop_exit/$exit
      -- CP-element group 64: 	 branch_block_stmt_546/do_while_stmt_547/loop_exit/ack
      -- 
    ack_864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_547_branch_ack_0, ack => writeEthernetHeaderToMem_CP_700_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	5 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_546/do_while_stmt_547/loop_taken/$exit
      -- CP-element group 65: 	 branch_block_stmt_546/do_while_stmt_547/loop_taken/ack
      -- 
    ack_868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_547_branch_ack_1, ack => writeEthernetHeaderToMem_CP_700_elements(65)); -- 
    -- CP-element group 66:  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	3 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	1 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_546/do_while_stmt_547/$exit
      -- 
    writeEthernetHeaderToMem_CP_700_elements(66) <= writeEthernetHeaderToMem_CP_700_elements(3);
    writeEthernetHeaderToMem_do_while_stmt_547_terminator_869: loop_terminator -- 
      generic map (name => " writeEthernetHeaderToMem_do_while_stmt_547_terminator_869", max_iterations_in_flight =>15) 
      port map(loop_body_exit => writeEthernetHeaderToMem_CP_700_elements(6),loop_continue => writeEthernetHeaderToMem_CP_700_elements(65),loop_terminate => writeEthernetHeaderToMem_CP_700_elements(64),loop_back => writeEthernetHeaderToMem_CP_700_elements(4),loop_exit => writeEthernetHeaderToMem_CP_700_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_549_phi_seq_783_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writeEthernetHeaderToMem_CP_700_elements(23);
      writeEthernetHeaderToMem_CP_700_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writeEthernetHeaderToMem_CP_700_elements(30);
      writeEthernetHeaderToMem_CP_700_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= writeEthernetHeaderToMem_CP_700_elements(31);
      writeEthernetHeaderToMem_CP_700_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= writeEthernetHeaderToMem_CP_700_elements(21);
      writeEthernetHeaderToMem_CP_700_elements(32)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writeEthernetHeaderToMem_CP_700_elements(34);
      writeEthernetHeaderToMem_CP_700_elements(33)<= src_update_reqs(1);
      src_update_acks(1)  <= writeEthernetHeaderToMem_CP_700_elements(35);
      writeEthernetHeaderToMem_CP_700_elements(22) <= phi_mux_reqs(1);
      phi_stmt_549_phi_seq_783 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_549_phi_seq_783") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writeEthernetHeaderToMem_CP_700_elements(17), 
          phi_sample_ack => writeEthernetHeaderToMem_CP_700_elements(18), 
          phi_update_req => writeEthernetHeaderToMem_CP_700_elements(19), 
          phi_update_ack => writeEthernetHeaderToMem_CP_700_elements(20), 
          phi_mux_ack => writeEthernetHeaderToMem_CP_700_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_555_phi_seq_827_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writeEthernetHeaderToMem_CP_700_elements(42);
      writeEthernetHeaderToMem_CP_700_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writeEthernetHeaderToMem_CP_700_elements(45);
      writeEthernetHeaderToMem_CP_700_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= writeEthernetHeaderToMem_CP_700_elements(47);
      writeEthernetHeaderToMem_CP_700_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= writeEthernetHeaderToMem_CP_700_elements(40);
      writeEthernetHeaderToMem_CP_700_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writeEthernetHeaderToMem_CP_700_elements(51);
      writeEthernetHeaderToMem_CP_700_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= writeEthernetHeaderToMem_CP_700_elements(52);
      writeEthernetHeaderToMem_CP_700_elements(41) <= phi_mux_reqs(1);
      phi_stmt_555_phi_seq_827 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_555_phi_seq_827") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writeEthernetHeaderToMem_CP_700_elements(11), 
          phi_sample_ack => writeEthernetHeaderToMem_CP_700_elements(38), 
          phi_update_req => writeEthernetHeaderToMem_CP_700_elements(13), 
          phi_update_ack => writeEthernetHeaderToMem_CP_700_elements(39), 
          phi_mux_ack => writeEthernetHeaderToMem_CP_700_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_725_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= writeEthernetHeaderToMem_CP_700_elements(7);
        preds(1)  <= writeEthernetHeaderToMem_CP_700_elements(8);
        entry_tmerge_725 : transition_merge -- 
          generic map(name => " entry_tmerge_725")
          port map (preds => preds, symbol_out => writeEthernetHeaderToMem_CP_700_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_553_wire : std_logic_vector(35 downto 0);
    signal I_555 : std_logic_vector(3 downto 0);
    signal RPIPE_nic_rx_to_header_562_wire : std_logic_vector(72 downto 0);
    signal ULE_u4_u1_597_wire : std_logic_vector(0 downto 0);
    signal ethernet_header_560 : std_logic_vector(72 downto 0);
    signal ignore_return_583 : std_logic_vector(63 downto 0);
    signal konst_552_wire_constant : std_logic_vector(35 downto 0);
    signal konst_586_wire_constant : std_logic_vector(3 downto 0);
    signal konst_591_wire_constant : std_logic_vector(35 downto 0);
    signal konst_596_wire_constant : std_logic_vector(3 downto 0);
    signal nI_588 : std_logic_vector(3 downto 0);
    signal nI_588_559_buffered : std_logic_vector(3 downto 0);
    signal nbuf_position_593 : std_logic_vector(35 downto 0);
    signal nbuf_position_593_554_buffered : std_logic_vector(35 downto 0);
    signal type_cast_558_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_576_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_578_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_570 : std_logic_vector(63 downto 0);
    signal wkeep_574 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_552_wire_constant <= "000000000000000000000000000000001000";
    konst_586_wire_constant <= "0001";
    konst_591_wire_constant <= "000000000000000000000000000000001000";
    konst_596_wire_constant <= "0001";
    type_cast_558_wire_constant <= "0000";
    type_cast_576_wire_constant <= "0";
    type_cast_578_wire_constant <= "0";
    phi_stmt_549: Block -- phi operator 
      signal idata: std_logic_vector(71 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u36_u36_553_wire & nbuf_position_593_554_buffered;
      req <= phi_stmt_549_req_0 & phi_stmt_549_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_549",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 36) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_549_ack_0,
          idata => idata,
          odata => buf_position_buffer,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_549
    phi_stmt_555: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_558_wire_constant & nI_588_559_buffered;
      req <= phi_stmt_555_req_0 & phi_stmt_555_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_555",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 4) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_555_ack_0,
          idata => idata,
          odata => I_555,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_555
    -- flow-through slice operator slice_569_inst
    wdata_570 <= ethernet_header_560(71 downto 8);
    -- flow-through slice operator slice_573_inst
    wkeep_574 <= ethernet_header_560(7 downto 0);
    nI_588_559_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nI_588_559_buf_req_0;
      nI_588_559_buf_ack_0<= wack(0);
      rreq(0) <= nI_588_559_buf_req_1;
      nI_588_559_buf_ack_1<= rack(0);
      nI_588_559_buf : InterlockBuffer generic map ( -- 
        name => "nI_588_559_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nI_588,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nI_588_559_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nbuf_position_593_554_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nbuf_position_593_554_buf_req_0;
      nbuf_position_593_554_buf_ack_0<= wack(0);
      rreq(0) <= nbuf_position_593_554_buf_req_1;
      nbuf_position_593_554_buf_ack_1<= rack(0);
      nbuf_position_593_554_buf : InterlockBuffer generic map ( -- 
        name => "nbuf_position_593_554_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nbuf_position_593,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nbuf_position_593_554_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_560
    process(RPIPE_nic_rx_to_header_562_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_nic_rx_to_header_562_wire(72 downto 0);
      ethernet_header_560 <= tmp_var; -- 
    end process;
    do_while_stmt_547_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULE_u4_u1_597_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_547_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_547_branch_req_0,
          ack0 => do_while_stmt_547_branch_ack_0,
          ack1 => do_while_stmt_547_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u36_u36_553_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= buf_pointer_buffer;
      ADD_u36_u36_553_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_553_inst_req_0;
      ADD_u36_u36_553_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_553_inst_req_1;
      ADD_u36_u36_553_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000001000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator ADD_u36_u36_592_inst
    process(buf_position_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buf_position_buffer, konst_591_wire_constant, tmp_var);
      nbuf_position_593 <= tmp_var; --
    end process;
    -- binary operator ADD_u4_u4_587_inst
    process(I_555) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApIntAdd_proc(I_555, konst_586_wire_constant, tmp_var);
      nI_588 <= tmp_var; --
    end process;
    -- binary operator ULE_u4_u1_597_inst
    process(nI_588) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(nI_588, konst_596_wire_constant, tmp_var);
      ULE_u4_u1_597_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_nic_rx_to_header_562_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_nic_rx_to_header_562_inst_req_0;
      RPIPE_nic_rx_to_header_562_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_nic_rx_to_header_562_inst_req_1;
      RPIPE_nic_rx_to_header_562_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_nic_rx_to_header_562_wire <= data_out(72 downto 0);
      nic_rx_to_header_read_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_header_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_header_read_0: InputPortRevised -- 
        generic map ( name => "nic_rx_to_header_read_0", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => nic_rx_to_header_pipe_read_req(0),
          oack => nic_rx_to_header_pipe_read_ack(0),
          odata => nic_rx_to_header_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared call operator group (0) : call_stmt_583_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 3);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_583_call_req_0;
      call_stmt_583_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_583_call_req_1;
      call_stmt_583_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_576_wire_constant & type_cast_578_wire_constant & wkeep_574 & buf_position_buffer & wdata_570;
      ignore_return_583 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writeEthernetHeaderToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity writePayloadToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    base_buf_pointer : in  std_logic_vector(35 downto 0);
    buf_pointer : in  std_logic_vector(35 downto 0);
    packet_size_32 : out  std_logic_vector(7 downto 0);
    bad_packet_identifier : out  std_logic_vector(0 downto 0);
    last_keep : out  std_logic_vector(7 downto 0);
    nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writePayloadToMem;
architecture writePayloadToMem_arch of writePayloadToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 72)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 17)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal base_buf_pointer_buffer :  std_logic_vector(35 downto 0);
  signal base_buf_pointer_update_enable: Boolean;
  signal buf_pointer_buffer :  std_logic_vector(35 downto 0);
  signal buf_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal packet_size_32_buffer :  std_logic_vector(7 downto 0);
  signal packet_size_32_update_enable: Boolean;
  signal bad_packet_identifier_buffer :  std_logic_vector(0 downto 0);
  signal bad_packet_identifier_update_enable: Boolean;
  signal last_keep_buffer :  std_logic_vector(7 downto 0);
  signal last_keep_update_enable: Boolean;
  signal writePayloadToMem_CP_870_start: Boolean;
  signal writePayloadToMem_CP_870_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_646_call_ack_0 : boolean;
  signal ADD_u36_u36_613_inst_req_1 : boolean;
  signal ADD_u36_u36_616_inst_req_0 : boolean;
  signal ADD_u36_u36_613_inst_ack_1 : boolean;
  signal phi_stmt_609_ack_0 : boolean;
  signal phi_stmt_609_req_1 : boolean;
  signal do_while_stmt_607_branch_req_0 : boolean;
  signal call_stmt_646_call_req_0 : boolean;
  signal RPIPE_nic_rx_to_packet_619_inst_ack_1 : boolean;
  signal ADD_u36_u36_613_inst_ack_0 : boolean;
  signal phi_stmt_609_req_0 : boolean;
  signal call_stmt_646_call_req_1 : boolean;
  signal RPIPE_nic_rx_to_packet_619_inst_req_1 : boolean;
  signal RPIPE_nic_rx_to_packet_619_inst_ack_0 : boolean;
  signal ADD_u36_u36_613_inst_req_0 : boolean;
  signal RPIPE_nic_rx_to_packet_619_inst_req_0 : boolean;
  signal do_while_stmt_607_branch_ack_1 : boolean;
  signal ADD_u36_u36_616_inst_ack_1 : boolean;
  signal do_while_stmt_607_branch_ack_0 : boolean;
  signal ADD_u36_u36_616_inst_req_1 : boolean;
  signal ADD_u36_u36_616_inst_ack_0 : boolean;
  signal call_stmt_646_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writePayloadToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 72) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= base_buf_pointer;
  base_buf_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(71 downto 36) <= buf_pointer;
  buf_pointer_buffer <= in_buffer_data_out(71 downto 36);
  in_buffer_data_in(tag_length + 71 downto 72) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 71 downto 72);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writePayloadToMem_CP_870_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writePayloadToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 17) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= packet_size_32_buffer;
  packet_size_32 <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(8 downto 8) <= bad_packet_identifier_buffer;
  bad_packet_identifier <= out_buffer_data_out(8 downto 8);
  out_buffer_data_in(16 downto 9) <= last_keep_buffer;
  last_keep <= out_buffer_data_out(16 downto 9);
  out_buffer_data_in(tag_length + 16 downto 17) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 16 downto 17);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writePayloadToMem_CP_870_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writePayloadToMem_CP_870_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writePayloadToMem_CP_870_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writePayloadToMem_CP_870: Block -- control-path 
    signal writePayloadToMem_CP_870_elements: BooleanArray(49 downto 0);
    -- 
  begin -- 
    writePayloadToMem_CP_870_elements(0) <= writePayloadToMem_CP_870_start;
    writePayloadToMem_CP_870_symbol <= writePayloadToMem_CP_870_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_606/do_while_stmt_607__entry__
      -- CP-element group 0: 	 branch_block_stmt_606/$entry
      -- CP-element group 0: 	 branch_block_stmt_606/branch_block_stmt_606__entry__
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	49 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_659_to_assign_stmt_674/$exit
      -- CP-element group 1: 	 assign_stmt_659_to_assign_stmt_674/$entry
      -- CP-element group 1: 	 branch_block_stmt_606/$exit
      -- CP-element group 1: 	 branch_block_stmt_606/do_while_stmt_607__exit__
      -- CP-element group 1: 	 branch_block_stmt_606/branch_block_stmt_606__exit__
      -- CP-element group 1: 	 $exit
      -- 
    writePayloadToMem_CP_870_elements(1) <= writePayloadToMem_CP_870_elements(49);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_606/do_while_stmt_607/$entry
      -- CP-element group 2: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607__entry__
      -- 
    writePayloadToMem_CP_870_elements(2) <= writePayloadToMem_CP_870_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	49 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607__exit__
      -- 
    -- Element group writePayloadToMem_CP_870_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_606/do_while_stmt_607/loop_back
      -- 
    -- Element group writePayloadToMem_CP_870_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	48 
    -- CP-element group 5: 	47 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_606/do_while_stmt_607/condition_done
      -- CP-element group 5: 	 branch_block_stmt_606/do_while_stmt_607/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_606/do_while_stmt_607/loop_exit/$entry
      -- 
    writePayloadToMem_CP_870_elements(5) <= writePayloadToMem_CP_870_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	46 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_606/do_while_stmt_607/loop_body_done
      -- 
    writePayloadToMem_CP_870_elements(6) <= writePayloadToMem_CP_870_elements(46);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/back_edge_to_loop_body
      -- 
    writePayloadToMem_CP_870_elements(7) <= writePayloadToMem_CP_870_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/first_time_through_loop_body
      -- 
    writePayloadToMem_CP_870_elements(8) <= writePayloadToMem_CP_870_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	36 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	45 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_617_sample_start_
      -- 
    -- Element group writePayloadToMem_CP_870_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	45 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/condition_evaluated
      -- 
    condition_evaluated_894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_870_elements(10), ack => do_while_stmt_607_branch_req_0); -- 
    writePayloadToMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_870_elements(14) & writePayloadToMem_CP_870_elements(45);
      gj_writePayloadToMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_870_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	37 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_609_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/aggregated_phi_sample_req
      -- 
    writePayloadToMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writePayloadToMem_CP_870_elements(9) & writePayloadToMem_CP_870_elements(15) & writePayloadToMem_CP_870_elements(14);
      gj_writePayloadToMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_870_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	39 
    -- CP-element group 12: 	17 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	46 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_609_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_617_sample_completed_
      -- 
    writePayloadToMem_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_870_elements(39) & writePayloadToMem_CP_870_elements(17);
      gj_writePayloadToMem_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_870_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	36 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	38 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_609_update_start__ps
      -- 
    writePayloadToMem_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_870_elements(36) & writePayloadToMem_CP_870_elements(16);
      gj_writePayloadToMem_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_870_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	40 
    -- CP-element group 14: 	18 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/aggregated_phi_update_ack
      -- 
    writePayloadToMem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_870_elements(40) & writePayloadToMem_CP_870_elements(18);
      gj_writePayloadToMem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_870_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_609_sample_start_
      -- 
    writePayloadToMem_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_870_elements(9) & writePayloadToMem_CP_870_elements(12);
      gj_writePayloadToMem_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_870_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	43 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_609_update_start_
      -- 
    writePayloadToMem_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_870_elements(9) & writePayloadToMem_CP_870_elements(43);
      gj_writePayloadToMem_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_870_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_609_sample_completed__ps
      -- 
    -- Element group writePayloadToMem_CP_870_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_609_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_609_update_completed__ps
      -- 
    -- Element group writePayloadToMem_CP_870_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_609_loopback_trigger
      -- 
    writePayloadToMem_CP_870_elements(19) <= writePayloadToMem_CP_870_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_609_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_609_loopback_sample_req_ps
      -- 
    phi_stmt_609_loopback_sample_req_909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_609_loopback_sample_req_909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_870_elements(20), ack => phi_stmt_609_req_1); -- 
    -- Element group writePayloadToMem_CP_870_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_609_entry_trigger
      -- 
    writePayloadToMem_CP_870_elements(21) <= writePayloadToMem_CP_870_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_609_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_609_entry_sample_req_ps
      -- 
    phi_stmt_609_entry_sample_req_912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_609_entry_sample_req_912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_870_elements(22), ack => phi_stmt_609_req_0); -- 
    -- Element group writePayloadToMem_CP_870_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_609_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_609_phi_mux_ack_ps
      -- 
    phi_stmt_609_phi_mux_ack_915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_609_ack_0, ack => writePayloadToMem_CP_870_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_613_sample_start__ps
      -- 
    -- Element group writePayloadToMem_CP_870_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_613_update_start__ps
      -- 
    -- Element group writePayloadToMem_CP_870_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_613_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_613_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_613_Sample/rr
      -- 
    rr_928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_870_elements(26), ack => ADD_u36_u36_613_inst_req_0); -- 
    writePayloadToMem_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_870_elements(24) & writePayloadToMem_CP_870_elements(28);
      gj_writePayloadToMem_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_870_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_613_Update/cr
      -- CP-element group 27: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_613_update_start_
      -- CP-element group 27: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_613_Update/$entry
      -- 
    cr_933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_870_elements(27), ack => ADD_u36_u36_613_inst_req_1); -- 
    writePayloadToMem_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_870_elements(25) & writePayloadToMem_CP_870_elements(29);
      gj_writePayloadToMem_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_870_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	26 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_613_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_613_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_613_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_613_Sample/$exit
      -- 
    ra_929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_613_inst_ack_0, ack => writePayloadToMem_CP_870_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_613_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_613_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_613_update_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_613_Update/$exit
      -- 
    ca_934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_613_inst_ack_1, ack => writePayloadToMem_CP_870_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_616_sample_start__ps
      -- 
    -- Element group writePayloadToMem_CP_870_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_616_update_start__ps
      -- 
    -- Element group writePayloadToMem_CP_870_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_616_Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_616_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_616_sample_start_
      -- 
    rr_946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_870_elements(32), ack => ADD_u36_u36_616_inst_req_0); -- 
    writePayloadToMem_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_870_elements(30) & writePayloadToMem_CP_870_elements(34);
      gj_writePayloadToMem_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_870_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	35 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_616_update_start_
      -- CP-element group 33: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_616_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_616_Update/$entry
      -- 
    cr_951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_870_elements(33), ack => ADD_u36_u36_616_inst_req_1); -- 
    writePayloadToMem_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_870_elements(31) & writePayloadToMem_CP_870_elements(35);
      gj_writePayloadToMem_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_870_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_616_sample_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_616_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_616_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_616_Sample/ra
      -- 
    ra_947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_616_inst_ack_0, ack => writePayloadToMem_CP_870_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	33 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_616_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_616_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_616_update_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/ADD_u36_u36_616_Update/$exit
      -- 
    ca_952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_616_inst_ack_1, ack => writePayloadToMem_CP_870_elements(35)); -- 
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	9 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	43 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	13 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_617_update_start_
      -- 
    writePayloadToMem_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_870_elements(9) & writePayloadToMem_CP_870_elements(43);
      gj_writePayloadToMem_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_870_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	11 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	40 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/RPIPE_nic_rx_to_packet_619_Sample/rr
      -- CP-element group 37: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/RPIPE_nic_rx_to_packet_619_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/RPIPE_nic_rx_to_packet_619_sample_start_
      -- 
    rr_965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_870_elements(37), ack => RPIPE_nic_rx_to_packet_619_inst_req_0); -- 
    writePayloadToMem_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_870_elements(11) & writePayloadToMem_CP_870_elements(40);
      gj_writePayloadToMem_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_870_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/RPIPE_nic_rx_to_packet_619_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/RPIPE_nic_rx_to_packet_619_Update/cr
      -- CP-element group 38: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/RPIPE_nic_rx_to_packet_619_update_start_
      -- 
    cr_970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_870_elements(38), ack => RPIPE_nic_rx_to_packet_619_inst_req_1); -- 
    writePayloadToMem_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_870_elements(39) & writePayloadToMem_CP_870_elements(13);
      gj_writePayloadToMem_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_870_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: 	12 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/RPIPE_nic_rx_to_packet_619_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/RPIPE_nic_rx_to_packet_619_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/RPIPE_nic_rx_to_packet_619_sample_completed_
      -- 
    ra_966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_packet_619_inst_ack_0, ack => writePayloadToMem_CP_870_elements(39)); -- 
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40: 	14 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	37 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/RPIPE_nic_rx_to_packet_619_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/RPIPE_nic_rx_to_packet_619_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/RPIPE_nic_rx_to_packet_619_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/phi_stmt_617_update_completed_
      -- 
    ca_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_packet_619_inst_ack_1, ack => writePayloadToMem_CP_870_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: 	18 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/call_stmt_646_Sample/crr
      -- CP-element group 41: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/call_stmt_646_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/call_stmt_646_sample_start_
      -- 
    crr_979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_870_elements(41), ack => call_stmt_646_call_req_0); -- 
    writePayloadToMem_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writePayloadToMem_CP_870_elements(40) & writePayloadToMem_CP_870_elements(18) & writePayloadToMem_CP_870_elements(43);
      gj_writePayloadToMem_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_870_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/call_stmt_646_update_start_
      -- CP-element group 42: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/call_stmt_646_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/call_stmt_646_Update/ccr
      -- 
    ccr_984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_870_elements(42), ack => call_stmt_646_call_req_1); -- 
    writePayloadToMem_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writePayloadToMem_CP_870_elements(44);
      gj_writePayloadToMem_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_870_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	41 
    -- CP-element group 43: 	16 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/call_stmt_646_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/call_stmt_646_Sample/cra
      -- CP-element group 43: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/call_stmt_646_Sample/$exit
      -- 
    cra_980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_646_call_ack_0, ack => writePayloadToMem_CP_870_elements(43)); -- 
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/call_stmt_646_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/call_stmt_646_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/call_stmt_646_Update/cca
      -- 
    cca_985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_646_call_ack_1, ack => writePayloadToMem_CP_870_elements(44)); -- 
    -- CP-element group 45:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	9 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	10 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group writePayloadToMem_CP_870_elements(45) is a control-delay.
    cp_element_45_delay: control_delay_element  generic map(name => " 45_delay", delay_value => 1)  port map(req => writePayloadToMem_CP_870_elements(9), ack => writePayloadToMem_CP_870_elements(45), clk => clk, reset =>reset);
    -- CP-element group 46:  join  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	12 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	6 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_606/do_while_stmt_607/do_while_stmt_607_loop_body/$exit
      -- 
    writePayloadToMem_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_870_elements(12) & writePayloadToMem_CP_870_elements(44);
      gj_writePayloadToMem_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_870_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	5 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_606/do_while_stmt_607/loop_exit/ack
      -- CP-element group 47: 	 branch_block_stmt_606/do_while_stmt_607/loop_exit/$exit
      -- 
    ack_990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_607_branch_ack_0, ack => writePayloadToMem_CP_870_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	5 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_606/do_while_stmt_607/loop_taken/ack
      -- CP-element group 48: 	 branch_block_stmt_606/do_while_stmt_607/loop_taken/$exit
      -- 
    ack_994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_607_branch_ack_1, ack => writePayloadToMem_CP_870_elements(48)); -- 
    -- CP-element group 49:  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	3 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	1 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_606/do_while_stmt_607/$exit
      -- 
    writePayloadToMem_CP_870_elements(49) <= writePayloadToMem_CP_870_elements(3);
    writePayloadToMem_do_while_stmt_607_terminator_995: loop_terminator -- 
      generic map (name => " writePayloadToMem_do_while_stmt_607_terminator_995", max_iterations_in_flight =>15) 
      port map(loop_body_exit => writePayloadToMem_CP_870_elements(6),loop_continue => writePayloadToMem_CP_870_elements(48),loop_terminate => writePayloadToMem_CP_870_elements(47),loop_back => writePayloadToMem_CP_870_elements(4),loop_exit => writePayloadToMem_CP_870_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_609_phi_seq_953_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writePayloadToMem_CP_870_elements(21);
      writePayloadToMem_CP_870_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writePayloadToMem_CP_870_elements(28);
      writePayloadToMem_CP_870_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= writePayloadToMem_CP_870_elements(29);
      writePayloadToMem_CP_870_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= writePayloadToMem_CP_870_elements(19);
      writePayloadToMem_CP_870_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writePayloadToMem_CP_870_elements(34);
      writePayloadToMem_CP_870_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= writePayloadToMem_CP_870_elements(35);
      writePayloadToMem_CP_870_elements(20) <= phi_mux_reqs(1);
      phi_stmt_609_phi_seq_953 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_609_phi_seq_953") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writePayloadToMem_CP_870_elements(11), 
          phi_sample_ack => writePayloadToMem_CP_870_elements(17), 
          phi_update_req => writePayloadToMem_CP_870_elements(13), 
          phi_update_ack => writePayloadToMem_CP_870_elements(18), 
          phi_mux_ack => writePayloadToMem_CP_870_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_895_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= writePayloadToMem_CP_870_elements(7);
        preds(1)  <= writePayloadToMem_CP_870_elements(8);
        entry_tmerge_895 : transition_merge -- 
          generic map(name => " entry_tmerge_895")
          port map (preds => preds, symbol_out => writePayloadToMem_CP_870_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_613_wire : std_logic_vector(35 downto 0);
    signal ADD_u36_u36_616_wire : std_logic_vector(35 downto 0);
    signal EQ_u64_u1_654_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_657_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_649_wire : std_logic_vector(0 downto 0);
    signal RPIPE_nic_rx_to_packet_619_wire : std_logic_vector(72 downto 0);
    signal R_BAD_PACKET_DATA_653_wire_constant : std_logic_vector(63 downto 0);
    signal SUB_u36_u36_663_wire : std_logic_vector(35 downto 0);
    signal buf_position_609 : std_logic_vector(35 downto 0);
    signal ignore_return_646 : std_logic_vector(63 downto 0);
    signal konst_612_wire_constant : std_logic_vector(35 downto 0);
    signal konst_615_wire_constant : std_logic_vector(35 downto 0);
    signal konst_656_wire_constant : std_logic_vector(7 downto 0);
    signal last_bit_624 : std_logic_vector(0 downto 0);
    signal packet_size_8_665 : std_logic_vector(7 downto 0);
    signal payload_data_617 : std_logic_vector(72 downto 0);
    signal type_cast_639_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_641_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_628 : std_logic_vector(63 downto 0);
    signal wkeep_632 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_BAD_PACKET_DATA_653_wire_constant <= "1111111111111111111111111111111111111111111111111111111111111111";
    konst_612_wire_constant <= "000000000000000000000000000000001000";
    konst_615_wire_constant <= "000000000000000000000000000000001000";
    konst_656_wire_constant <= "00000000";
    type_cast_639_wire_constant <= "0";
    type_cast_641_wire_constant <= "0";
    phi_stmt_609: Block -- phi operator 
      signal idata: std_logic_vector(71 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u36_u36_613_wire & ADD_u36_u36_616_wire;
      req <= phi_stmt_609_req_0 & phi_stmt_609_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_609",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 36) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_609_ack_0,
          idata => idata,
          odata => buf_position_609,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_609
    -- flow-through slice operator slice_623_inst
    last_bit_624 <= payload_data_617(72 downto 72);
    -- flow-through slice operator slice_627_inst
    wdata_628 <= payload_data_617(71 downto 8);
    -- flow-through slice operator slice_631_inst
    wkeep_632 <= payload_data_617(7 downto 0);
    -- interlock W_last_keep_672_inst
    process(wkeep_632) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := wkeep_632(7 downto 0);
      last_keep_buffer <= tmp_var; -- 
    end process;
    -- interlock W_packet_size_32_666_inst
    process(packet_size_8_665) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := packet_size_8_665(7 downto 0);
      packet_size_32_buffer <= tmp_var; -- 
    end process;
    -- interlock ssrc_phi_stmt_617
    process(RPIPE_nic_rx_to_packet_619_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_nic_rx_to_packet_619_wire(72 downto 0);
      payload_data_617 <= tmp_var; -- 
    end process;
    -- interlock type_cast_664_inst
    process(SUB_u36_u36_663_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := SUB_u36_u36_663_wire(7 downto 0);
      packet_size_8_665 <= tmp_var; -- 
    end process;
    do_while_stmt_607_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_649_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_607_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_607_branch_req_0,
          ack0 => do_while_stmt_607_branch_ack_0,
          ack1 => do_while_stmt_607_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u36_u36_613_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= buf_pointer_buffer;
      ADD_u36_u36_613_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_613_inst_req_0;
      ADD_u36_u36_613_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_613_inst_req_1;
      ADD_u36_u36_613_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000001000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : ADD_u36_u36_616_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= buf_position_609;
      ADD_u36_u36_616_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_616_inst_req_0;
      ADD_u36_u36_616_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_616_inst_req_1;
      ADD_u36_u36_616_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000001000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- binary operator AND_u1_u1_658_inst
    process(EQ_u64_u1_654_wire, EQ_u8_u1_657_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u64_u1_654_wire, EQ_u8_u1_657_wire, tmp_var);
      bad_packet_identifier_buffer <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_654_inst
    process(wdata_628) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(wdata_628, R_BAD_PACKET_DATA_653_wire_constant, tmp_var);
      EQ_u64_u1_654_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_657_inst
    process(wkeep_632) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(wkeep_632, konst_656_wire_constant, tmp_var);
      EQ_u8_u1_657_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_649_inst
    process(last_bit_624) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", last_bit_624, tmp_var);
      NOT_u1_u1_649_wire <= tmp_var; -- 
    end process;
    -- binary operator SUB_u36_u36_663_inst
    process(buf_position_609, base_buf_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntSub_proc(buf_position_609, base_buf_pointer_buffer, tmp_var);
      SUB_u36_u36_663_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_nic_rx_to_packet_619_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_nic_rx_to_packet_619_inst_req_0;
      RPIPE_nic_rx_to_packet_619_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_nic_rx_to_packet_619_inst_req_1;
      RPIPE_nic_rx_to_packet_619_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_nic_rx_to_packet_619_wire <= data_out(72 downto 0);
      nic_rx_to_packet_read_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_packet_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_packet_read_0: InputPortRevised -- 
        generic map ( name => "nic_rx_to_packet_read_0", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => nic_rx_to_packet_pipe_read_req(0),
          oack => nic_rx_to_packet_pipe_read_ack(0),
          odata => nic_rx_to_packet_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared call operator group (0) : call_stmt_646_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 3);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_646_call_req_0;
      call_stmt_646_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_646_call_req_1;
      call_stmt_646_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_639_wire_constant & type_cast_641_wire_constant & wkeep_632 & buf_position_609 & wdata_628;
      ignore_return_646 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writePayloadToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    AFB_NIC_REQUEST_pipe_write_data: in std_logic_vector(73 downto 0);
    AFB_NIC_REQUEST_pipe_write_req : in std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_write_ack : out std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_read_data: out std_logic_vector(32 downto 0);
    AFB_NIC_RESPONSE_pipe_read_req : in std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_read_ack : out std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_data: in std_logic_vector(64 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_req : in std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_ack : out std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_data: out std_logic_vector(109 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_req : in std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_ack : out std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_write_data: in std_logic_vector(72 downto 0);
    mac_to_nic_data_pipe_write_req : in std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_write_ack : out std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_data: out std_logic_vector(72 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(11 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(39 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(5 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(5 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(2 downto 0);
  -- declarations related to module AccessRegister
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module AccessRegister
  signal AccessRegister_rwbar :  std_logic_vector(0 downto 0);
  signal AccessRegister_bmask :  std_logic_vector(3 downto 0);
  signal AccessRegister_register_index :  std_logic_vector(5 downto 0);
  signal AccessRegister_wdata :  std_logic_vector(31 downto 0);
  signal AccessRegister_rdata :  std_logic_vector(31 downto 0);
  signal AccessRegister_in_args    : std_logic_vector(42 downto 0);
  signal AccessRegister_out_args   : std_logic_vector(31 downto 0);
  signal AccessRegister_tag_in    : std_logic_vector(4 downto 0) := (others => '0');
  signal AccessRegister_tag_out   : std_logic_vector(4 downto 0);
  signal AccessRegister_start_req : std_logic;
  signal AccessRegister_start_ack : std_logic;
  signal AccessRegister_fin_req   : std_logic;
  signal AccessRegister_fin_ack : std_logic;
  -- caller side aggregated signals for module AccessRegister
  signal AccessRegister_call_reqs: std_logic_vector(3 downto 0);
  signal AccessRegister_call_acks: std_logic_vector(3 downto 0);
  signal AccessRegister_return_reqs: std_logic_vector(3 downto 0);
  signal AccessRegister_return_acks: std_logic_vector(3 downto 0);
  signal AccessRegister_call_data: std_logic_vector(171 downto 0);
  signal AccessRegister_call_tag: std_logic_vector(7 downto 0);
  signal AccessRegister_return_data: std_logic_vector(127 downto 0);
  signal AccessRegister_return_tag: std_logic_vector(7 downto 0);
  -- declarations related to module NicRegisterAccessDaemon
  component NicRegisterAccessDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(42 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(32 downto 0);
      UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
      UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
      UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module NicRegisterAccessDaemon
  signal NicRegisterAccessDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal NicRegisterAccessDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal NicRegisterAccessDaemon_start_req : std_logic;
  signal NicRegisterAccessDaemon_start_ack : std_logic;
  signal NicRegisterAccessDaemon_fin_req   : std_logic;
  signal NicRegisterAccessDaemon_fin_ack : std_logic;
  -- declarations related to module ReceiveEngineDaemon
  component ReceiveEngineDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      FREE_Q : in std_logic_vector(35 downto 0);
      CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
      populateRxQueue_call_reqs : out  std_logic_vector(0 downto 0);
      populateRxQueue_call_acks : in   std_logic_vector(0 downto 0);
      populateRxQueue_call_data : out  std_logic_vector(35 downto 0);
      populateRxQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      populateRxQueue_return_reqs : out  std_logic_vector(0 downto 0);
      populateRxQueue_return_acks : in   std_logic_vector(0 downto 0);
      populateRxQueue_return_tag :  in   std_logic_vector(0 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(36 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(32 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      loadBuffer_call_reqs : out  std_logic_vector(0 downto 0);
      loadBuffer_call_acks : in   std_logic_vector(0 downto 0);
      loadBuffer_call_data : out  std_logic_vector(35 downto 0);
      loadBuffer_call_tag  :  out  std_logic_vector(0 downto 0);
      loadBuffer_return_reqs : out  std_logic_vector(0 downto 0);
      loadBuffer_return_acks : in   std_logic_vector(0 downto 0);
      loadBuffer_return_data : in   std_logic_vector(0 downto 0);
      loadBuffer_return_tag :  in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module ReceiveEngineDaemon
  signal ReceiveEngineDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal ReceiveEngineDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal ReceiveEngineDaemon_start_req : std_logic;
  signal ReceiveEngineDaemon_start_ack : std_logic;
  signal ReceiveEngineDaemon_fin_req   : std_logic;
  signal ReceiveEngineDaemon_fin_ack : std_logic;
  -- declarations related to module SoftwareRegisterAccessDaemon
  component SoftwareRegisterAccessDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      AFB_NIC_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
      AFB_NIC_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
      AFB_NIC_REQUEST_pipe_read_data : in   std_logic_vector(73 downto 0);
      FREE_Q_pipe_write_req : out  std_logic_vector(0 downto 0);
      FREE_Q_pipe_write_ack : in   std_logic_vector(0 downto 0);
      FREE_Q_pipe_write_data : out  std_logic_vector(35 downto 0);
      AFB_NIC_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
      AFB_NIC_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      AFB_NIC_RESPONSE_pipe_write_data : out  std_logic_vector(32 downto 0);
      CONTROL_REGISTER_pipe_write_req : out  std_logic_vector(0 downto 0);
      CONTROL_REGISTER_pipe_write_ack : in   std_logic_vector(0 downto 0);
      CONTROL_REGISTER_pipe_write_data : out  std_logic_vector(31 downto 0);
      NUMBER_OF_SERVERS_pipe_write_req : out  std_logic_vector(0 downto 0);
      NUMBER_OF_SERVERS_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NUMBER_OF_SERVERS_pipe_write_data : out  std_logic_vector(31 downto 0);
      UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
      UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
      UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module SoftwareRegisterAccessDaemon
  signal SoftwareRegisterAccessDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal SoftwareRegisterAccessDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal SoftwareRegisterAccessDaemon_start_req : std_logic;
  signal SoftwareRegisterAccessDaemon_start_ack : std_logic;
  signal SoftwareRegisterAccessDaemon_fin_req   : std_logic;
  signal SoftwareRegisterAccessDaemon_fin_ack : std_logic;
  -- declarations related to module UpdateRegister
  component UpdateRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      bmask : in  std_logic_vector(3 downto 0);
      rval : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      index : in  std_logic_vector(5 downto 0);
      wval : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module UpdateRegister
  signal UpdateRegister_bmask :  std_logic_vector(3 downto 0);
  signal UpdateRegister_rval :  std_logic_vector(31 downto 0);
  signal UpdateRegister_wdata :  std_logic_vector(31 downto 0);
  signal UpdateRegister_index :  std_logic_vector(5 downto 0);
  signal UpdateRegister_wval :  std_logic_vector(31 downto 0);
  signal UpdateRegister_in_args    : std_logic_vector(73 downto 0);
  signal UpdateRegister_out_args   : std_logic_vector(31 downto 0);
  signal UpdateRegister_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal UpdateRegister_tag_out   : std_logic_vector(2 downto 0);
  signal UpdateRegister_start_req : std_logic;
  signal UpdateRegister_start_ack : std_logic;
  signal UpdateRegister_fin_req   : std_logic;
  signal UpdateRegister_fin_ack : std_logic;
  -- caller side aggregated signals for module UpdateRegister
  signal UpdateRegister_call_reqs: std_logic_vector(1 downto 0);
  signal UpdateRegister_call_acks: std_logic_vector(1 downto 0);
  signal UpdateRegister_return_reqs: std_logic_vector(1 downto 0);
  signal UpdateRegister_return_acks: std_logic_vector(1 downto 0);
  signal UpdateRegister_call_data: std_logic_vector(147 downto 0);
  signal UpdateRegister_call_tag: std_logic_vector(1 downto 0);
  signal UpdateRegister_return_data: std_logic_vector(63 downto 0);
  signal UpdateRegister_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module accessMemory
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMemory
  signal accessMemory_lock :  std_logic_vector(0 downto 0);
  signal accessMemory_rwbar :  std_logic_vector(0 downto 0);
  signal accessMemory_bmask :  std_logic_vector(7 downto 0);
  signal accessMemory_addr :  std_logic_vector(35 downto 0);
  signal accessMemory_wdata :  std_logic_vector(63 downto 0);
  signal accessMemory_rdata :  std_logic_vector(63 downto 0);
  signal accessMemory_in_args    : std_logic_vector(109 downto 0);
  signal accessMemory_out_args   : std_logic_vector(63 downto 0);
  signal accessMemory_tag_in    : std_logic_vector(5 downto 0) := (others => '0');
  signal accessMemory_tag_out   : std_logic_vector(5 downto 0);
  signal accessMemory_start_req : std_logic;
  signal accessMemory_start_ack : std_logic;
  signal accessMemory_fin_req   : std_logic;
  signal accessMemory_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMemory
  signal accessMemory_call_reqs: std_logic_vector(10 downto 0);
  signal accessMemory_call_acks: std_logic_vector(10 downto 0);
  signal accessMemory_return_reqs: std_logic_vector(10 downto 0);
  signal accessMemory_return_acks: std_logic_vector(10 downto 0);
  signal accessMemory_call_data: std_logic_vector(1209 downto 0);
  signal accessMemory_call_tag: std_logic_vector(21 downto 0);
  signal accessMemory_return_data: std_logic_vector(703 downto 0);
  signal accessMemory_return_tag: std_logic_vector(21 downto 0);
  -- declarations related to module acquireMutex
  component acquireMutex is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module acquireMutex
  signal acquireMutex_q_base_address :  std_logic_vector(35 downto 0);
  signal acquireMutex_m_ok :  std_logic_vector(0 downto 0);
  signal acquireMutex_in_args    : std_logic_vector(35 downto 0);
  signal acquireMutex_out_args   : std_logic_vector(0 downto 0);
  signal acquireMutex_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal acquireMutex_tag_out   : std_logic_vector(2 downto 0);
  signal acquireMutex_start_req : std_logic;
  signal acquireMutex_start_ack : std_logic;
  signal acquireMutex_fin_req   : std_logic;
  signal acquireMutex_fin_ack : std_logic;
  -- caller side aggregated signals for module acquireMutex
  signal acquireMutex_call_reqs: std_logic_vector(1 downto 0);
  signal acquireMutex_call_acks: std_logic_vector(1 downto 0);
  signal acquireMutex_return_reqs: std_logic_vector(1 downto 0);
  signal acquireMutex_return_acks: std_logic_vector(1 downto 0);
  signal acquireMutex_call_data: std_logic_vector(71 downto 0);
  signal acquireMutex_call_tag: std_logic_vector(1 downto 0);
  signal acquireMutex_return_data: std_logic_vector(1 downto 0);
  signal acquireMutex_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module delay_time
  -- declarations related to module getQueueElement
  component getQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      read_pointer : in  std_logic_vector(31 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueueElement
  signal getQueueElement_q_base_address :  std_logic_vector(35 downto 0);
  signal getQueueElement_read_pointer :  std_logic_vector(31 downto 0);
  signal getQueueElement_q_r_data :  std_logic_vector(31 downto 0);
  signal getQueueElement_in_args    : std_logic_vector(67 downto 0);
  signal getQueueElement_out_args   : std_logic_vector(31 downto 0);
  signal getQueueElement_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal getQueueElement_tag_out   : std_logic_vector(1 downto 0);
  signal getQueueElement_start_req : std_logic;
  signal getQueueElement_start_ack : std_logic;
  signal getQueueElement_fin_req   : std_logic;
  signal getQueueElement_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueueElement
  signal getQueueElement_call_reqs: std_logic_vector(0 downto 0);
  signal getQueueElement_call_acks: std_logic_vector(0 downto 0);
  signal getQueueElement_return_reqs: std_logic_vector(0 downto 0);
  signal getQueueElement_return_acks: std_logic_vector(0 downto 0);
  signal getQueueElement_call_data: std_logic_vector(67 downto 0);
  signal getQueueElement_call_tag: std_logic_vector(0 downto 0);
  signal getQueueElement_return_data: std_logic_vector(31 downto 0);
  signal getQueueElement_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module getQueuePointers
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueuePointers
  signal getQueuePointers_q_base_address :  std_logic_vector(35 downto 0);
  signal getQueuePointers_wp :  std_logic_vector(31 downto 0);
  signal getQueuePointers_rp :  std_logic_vector(31 downto 0);
  signal getQueuePointers_in_args    : std_logic_vector(35 downto 0);
  signal getQueuePointers_out_args   : std_logic_vector(63 downto 0);
  signal getQueuePointers_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal getQueuePointers_tag_out   : std_logic_vector(2 downto 0);
  signal getQueuePointers_start_req : std_logic;
  signal getQueuePointers_start_ack : std_logic;
  signal getQueuePointers_fin_req   : std_logic;
  signal getQueuePointers_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueuePointers
  signal getQueuePointers_call_reqs: std_logic_vector(1 downto 0);
  signal getQueuePointers_call_acks: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_reqs: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_acks: std_logic_vector(1 downto 0);
  signal getQueuePointers_call_data: std_logic_vector(71 downto 0);
  signal getQueuePointers_call_tag: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_data: std_logic_vector(127 downto 0);
  signal getQueuePointers_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module getTxPacketPointerFromServer
  component getTxPacketPointerFromServer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_index : in  std_logic_vector(5 downto 0);
      pkt_pointer : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(36 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(32 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getTxPacketPointerFromServer
  signal getTxPacketPointerFromServer_queue_index :  std_logic_vector(5 downto 0);
  signal getTxPacketPointerFromServer_pkt_pointer :  std_logic_vector(31 downto 0);
  signal getTxPacketPointerFromServer_status :  std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_in_args    : std_logic_vector(5 downto 0);
  signal getTxPacketPointerFromServer_out_args   : std_logic_vector(32 downto 0);
  signal getTxPacketPointerFromServer_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal getTxPacketPointerFromServer_tag_out   : std_logic_vector(1 downto 0);
  signal getTxPacketPointerFromServer_start_req : std_logic;
  signal getTxPacketPointerFromServer_start_ack : std_logic;
  signal getTxPacketPointerFromServer_fin_req   : std_logic;
  signal getTxPacketPointerFromServer_fin_ack : std_logic;
  -- caller side aggregated signals for module getTxPacketPointerFromServer
  signal getTxPacketPointerFromServer_call_reqs: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_call_acks: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_reqs: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_acks: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_call_data: std_logic_vector(5 downto 0);
  signal getTxPacketPointerFromServer_call_tag: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_data: std_logic_vector(32 downto 0);
  signal getTxPacketPointerFromServer_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module loadBuffer
  component loadBuffer is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_data : out  std_logic_vector(51 downto 0);
      writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_data : out  std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_data : in   std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_data : out  std_logic_vector(71 downto 0);
      writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_return_data : in   std_logic_vector(16 downto 0);
      writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadBuffer
  signal loadBuffer_rx_buffer_pointer :  std_logic_vector(35 downto 0);
  signal loadBuffer_bad_packet_identifier :  std_logic_vector(0 downto 0);
  signal loadBuffer_in_args    : std_logic_vector(35 downto 0);
  signal loadBuffer_out_args   : std_logic_vector(0 downto 0);
  signal loadBuffer_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadBuffer_tag_out   : std_logic_vector(1 downto 0);
  signal loadBuffer_start_req : std_logic;
  signal loadBuffer_start_ack : std_logic;
  signal loadBuffer_fin_req   : std_logic;
  signal loadBuffer_fin_ack : std_logic;
  -- caller side aggregated signals for module loadBuffer
  signal loadBuffer_call_reqs: std_logic_vector(0 downto 0);
  signal loadBuffer_call_acks: std_logic_vector(0 downto 0);
  signal loadBuffer_return_reqs: std_logic_vector(0 downto 0);
  signal loadBuffer_return_acks: std_logic_vector(0 downto 0);
  signal loadBuffer_call_data: std_logic_vector(35 downto 0);
  signal loadBuffer_call_tag: std_logic_vector(0 downto 0);
  signal loadBuffer_return_data: std_logic_vector(0 downto 0);
  signal loadBuffer_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module nextLSTATE
  -- declarations related to module nicRxFromMacDaemon
  component nicRxFromMacDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      mac_to_nic_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      mac_to_nic_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      mac_to_nic_data_pipe_read_data : in   std_logic_vector(72 downto 0);
      CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      nic_rx_to_packet_pipe_write_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_write_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_write_data : out  std_logic_vector(72 downto 0);
      nic_rx_to_header_pipe_write_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_write_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_write_data : out  std_logic_vector(72 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module nicRxFromMacDaemon
  signal nicRxFromMacDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal nicRxFromMacDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal nicRxFromMacDaemon_start_req : std_logic;
  signal nicRxFromMacDaemon_start_ack : std_logic;
  signal nicRxFromMacDaemon_fin_req   : std_logic;
  signal nicRxFromMacDaemon_fin_ack : std_logic;
  -- declarations related to module popFromQueue
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(67 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(31 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module popFromQueue
  signal popFromQueue_lock :  std_logic_vector(0 downto 0);
  signal popFromQueue_q_base_address :  std_logic_vector(35 downto 0);
  signal popFromQueue_q_r_data :  std_logic_vector(31 downto 0);
  signal popFromQueue_status :  std_logic_vector(0 downto 0);
  signal popFromQueue_in_args    : std_logic_vector(36 downto 0);
  signal popFromQueue_out_args   : std_logic_vector(32 downto 0);
  signal popFromQueue_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal popFromQueue_tag_out   : std_logic_vector(2 downto 0);
  signal popFromQueue_start_req : std_logic;
  signal popFromQueue_start_ack : std_logic;
  signal popFromQueue_fin_req   : std_logic;
  signal popFromQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module popFromQueue
  signal popFromQueue_call_reqs: std_logic_vector(1 downto 0);
  signal popFromQueue_call_acks: std_logic_vector(1 downto 0);
  signal popFromQueue_return_reqs: std_logic_vector(1 downto 0);
  signal popFromQueue_return_acks: std_logic_vector(1 downto 0);
  signal popFromQueue_call_data: std_logic_vector(73 downto 0);
  signal popFromQueue_call_tag: std_logic_vector(1 downto 0);
  signal popFromQueue_return_data: std_logic_vector(65 downto 0);
  signal popFromQueue_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module populateRxQueue
  component populateRxQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
      NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module populateRxQueue
  signal populateRxQueue_rx_buffer_pointer :  std_logic_vector(35 downto 0);
  signal populateRxQueue_in_args    : std_logic_vector(35 downto 0);
  signal populateRxQueue_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal populateRxQueue_tag_out   : std_logic_vector(1 downto 0);
  signal populateRxQueue_start_req : std_logic;
  signal populateRxQueue_start_ack : std_logic;
  signal populateRxQueue_fin_req   : std_logic;
  signal populateRxQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module populateRxQueue
  signal populateRxQueue_call_reqs: std_logic_vector(0 downto 0);
  signal populateRxQueue_call_acks: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_reqs: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_acks: std_logic_vector(0 downto 0);
  signal populateRxQueue_call_data: std_logic_vector(35 downto 0);
  signal populateRxQueue_call_tag: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module pushIntoQueue
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module pushIntoQueue
  signal pushIntoQueue_lock :  std_logic_vector(0 downto 0);
  signal pushIntoQueue_q_base_address :  std_logic_vector(35 downto 0);
  signal pushIntoQueue_q_w_data :  std_logic_vector(31 downto 0);
  signal pushIntoQueue_status :  std_logic_vector(0 downto 0);
  signal pushIntoQueue_in_args    : std_logic_vector(68 downto 0);
  signal pushIntoQueue_out_args   : std_logic_vector(0 downto 0);
  signal pushIntoQueue_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal pushIntoQueue_tag_out   : std_logic_vector(2 downto 0);
  signal pushIntoQueue_start_req : std_logic;
  signal pushIntoQueue_start_ack : std_logic;
  signal pushIntoQueue_fin_req   : std_logic;
  signal pushIntoQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module pushIntoQueue
  signal pushIntoQueue_call_reqs: std_logic_vector(2 downto 0);
  signal pushIntoQueue_call_acks: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_reqs: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_acks: std_logic_vector(2 downto 0);
  signal pushIntoQueue_call_data: std_logic_vector(206 downto 0);
  signal pushIntoQueue_call_tag: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_data: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_tag: std_logic_vector(2 downto 0);
  -- declarations related to module releaseMutex
  component releaseMutex is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module releaseMutex
  signal releaseMutex_q_base_address :  std_logic_vector(35 downto 0);
  signal releaseMutex_in_args    : std_logic_vector(35 downto 0);
  signal releaseMutex_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal releaseMutex_tag_out   : std_logic_vector(2 downto 0);
  signal releaseMutex_start_req : std_logic;
  signal releaseMutex_start_ack : std_logic;
  signal releaseMutex_fin_req   : std_logic;
  signal releaseMutex_fin_ack : std_logic;
  -- caller side aggregated signals for module releaseMutex
  signal releaseMutex_call_reqs: std_logic_vector(1 downto 0);
  signal releaseMutex_call_acks: std_logic_vector(1 downto 0);
  signal releaseMutex_return_reqs: std_logic_vector(1 downto 0);
  signal releaseMutex_return_acks: std_logic_vector(1 downto 0);
  signal releaseMutex_call_data: std_logic_vector(71 downto 0);
  signal releaseMutex_call_tag: std_logic_vector(1 downto 0);
  signal releaseMutex_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module setQueueElement
  component setQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      write_pointer : in  std_logic_vector(31 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module setQueueElement
  signal setQueueElement_q_base_address :  std_logic_vector(35 downto 0);
  signal setQueueElement_write_pointer :  std_logic_vector(31 downto 0);
  signal setQueueElement_q_w_data :  std_logic_vector(31 downto 0);
  signal setQueueElement_in_args    : std_logic_vector(99 downto 0);
  signal setQueueElement_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal setQueueElement_tag_out   : std_logic_vector(1 downto 0);
  signal setQueueElement_start_req : std_logic;
  signal setQueueElement_start_ack : std_logic;
  signal setQueueElement_fin_req   : std_logic;
  signal setQueueElement_fin_ack : std_logic;
  -- caller side aggregated signals for module setQueueElement
  signal setQueueElement_call_reqs: std_logic_vector(0 downto 0);
  signal setQueueElement_call_acks: std_logic_vector(0 downto 0);
  signal setQueueElement_return_reqs: std_logic_vector(0 downto 0);
  signal setQueueElement_return_acks: std_logic_vector(0 downto 0);
  signal setQueueElement_call_data: std_logic_vector(99 downto 0);
  signal setQueueElement_call_tag: std_logic_vector(0 downto 0);
  signal setQueueElement_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module setQueuePointers
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module setQueuePointers
  signal setQueuePointers_q_base_address :  std_logic_vector(35 downto 0);
  signal setQueuePointers_wp :  std_logic_vector(31 downto 0);
  signal setQueuePointers_rp :  std_logic_vector(31 downto 0);
  signal setQueuePointers_in_args    : std_logic_vector(99 downto 0);
  signal setQueuePointers_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal setQueuePointers_tag_out   : std_logic_vector(2 downto 0);
  signal setQueuePointers_start_req : std_logic;
  signal setQueuePointers_start_ack : std_logic;
  signal setQueuePointers_fin_req   : std_logic;
  signal setQueuePointers_fin_ack : std_logic;
  -- caller side aggregated signals for module setQueuePointers
  signal setQueuePointers_call_reqs: std_logic_vector(1 downto 0);
  signal setQueuePointers_call_acks: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_reqs: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_acks: std_logic_vector(1 downto 0);
  signal setQueuePointers_call_data: std_logic_vector(199 downto 0);
  signal setQueuePointers_call_tag: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module transmitEngineDaemon
  component transmitEngineDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      FREE_Q : in std_logic_vector(35 downto 0);
      LAST_READ_TX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
      CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(1 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(1 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(11 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_reqs : out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_acks : in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_data : out  std_logic_vector(5 downto 0);
      getTxPacketPointerFromServer_call_tag  :  out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_reqs : out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_acks : in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_data : in   std_logic_vector(32 downto 0);
      getTxPacketPointerFromServer_return_tag :  in   std_logic_vector(0 downto 0);
      transmitPacket_call_reqs : out  std_logic_vector(0 downto 0);
      transmitPacket_call_acks : in   std_logic_vector(0 downto 0);
      transmitPacket_call_data : out  std_logic_vector(31 downto 0);
      transmitPacket_call_tag  :  out  std_logic_vector(0 downto 0);
      transmitPacket_return_reqs : out  std_logic_vector(0 downto 0);
      transmitPacket_return_acks : in   std_logic_vector(0 downto 0);
      transmitPacket_return_data : in   std_logic_vector(0 downto 0);
      transmitPacket_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module transmitEngineDaemon
  signal transmitEngineDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal transmitEngineDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal transmitEngineDaemon_start_req : std_logic;
  signal transmitEngineDaemon_start_ack : std_logic;
  signal transmitEngineDaemon_fin_req   : std_logic;
  signal transmitEngineDaemon_fin_ack : std_logic;
  -- declarations related to module transmitPacket
  component transmitPacket is -- 
    generic (tag_length : integer); 
    port ( -- 
      packet_pointer : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(145 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_call_acks : in   std_logic_vector(1 downto 0);
      accessMemory_call_data : out  std_logic_vector(219 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(3 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_return_acks : in   std_logic_vector(1 downto 0);
      accessMemory_return_data : in   std_logic_vector(127 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module transmitPacket
  signal transmitPacket_packet_pointer :  std_logic_vector(31 downto 0);
  signal transmitPacket_status :  std_logic_vector(0 downto 0);
  signal transmitPacket_in_args    : std_logic_vector(31 downto 0);
  signal transmitPacket_out_args   : std_logic_vector(0 downto 0);
  signal transmitPacket_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal transmitPacket_tag_out   : std_logic_vector(1 downto 0);
  signal transmitPacket_start_req : std_logic;
  signal transmitPacket_start_ack : std_logic;
  signal transmitPacket_fin_req   : std_logic;
  signal transmitPacket_fin_ack : std_logic;
  -- caller side aggregated signals for module transmitPacket
  signal transmitPacket_call_reqs: std_logic_vector(0 downto 0);
  signal transmitPacket_call_acks: std_logic_vector(0 downto 0);
  signal transmitPacket_return_reqs: std_logic_vector(0 downto 0);
  signal transmitPacket_return_acks: std_logic_vector(0 downto 0);
  signal transmitPacket_call_data: std_logic_vector(31 downto 0);
  signal transmitPacket_call_tag: std_logic_vector(0 downto 0);
  signal transmitPacket_return_data: std_logic_vector(0 downto 0);
  signal transmitPacket_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writeControlInformationToMem
  component writeControlInformationToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buffer_pointer : in  std_logic_vector(35 downto 0);
      packet_size : in  std_logic_vector(7 downto 0);
      last_keep : in  std_logic_vector(7 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeControlInformationToMem
  signal writeControlInformationToMem_base_buffer_pointer :  std_logic_vector(35 downto 0);
  signal writeControlInformationToMem_packet_size :  std_logic_vector(7 downto 0);
  signal writeControlInformationToMem_last_keep :  std_logic_vector(7 downto 0);
  signal writeControlInformationToMem_in_args    : std_logic_vector(51 downto 0);
  signal writeControlInformationToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeControlInformationToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writeControlInformationToMem_start_req : std_logic;
  signal writeControlInformationToMem_start_ack : std_logic;
  signal writeControlInformationToMem_fin_req   : std_logic;
  signal writeControlInformationToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writeControlInformationToMem
  signal writeControlInformationToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_call_acks: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_acks: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_call_data: std_logic_vector(51 downto 0);
  signal writeControlInformationToMem_call_tag: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writeEthernetHeaderToMem
  component writeEthernetHeaderToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      buf_pointer : in  std_logic_vector(35 downto 0);
      buf_position : out  std_logic_vector(35 downto 0);
      nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeEthernetHeaderToMem
  signal writeEthernetHeaderToMem_buf_pointer :  std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_buf_position :  std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_in_args    : std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_out_args   : std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeEthernetHeaderToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writeEthernetHeaderToMem_start_req : std_logic;
  signal writeEthernetHeaderToMem_start_ack : std_logic;
  signal writeEthernetHeaderToMem_fin_req   : std_logic;
  signal writeEthernetHeaderToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writeEthernetHeaderToMem
  signal writeEthernetHeaderToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_call_acks: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_acks: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_call_data: std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_call_tag: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_data: std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writePayloadToMem
  component writePayloadToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buf_pointer : in  std_logic_vector(35 downto 0);
      buf_pointer : in  std_logic_vector(35 downto 0);
      packet_size_32 : out  std_logic_vector(7 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      last_keep : out  std_logic_vector(7 downto 0);
      nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writePayloadToMem
  signal writePayloadToMem_base_buf_pointer :  std_logic_vector(35 downto 0);
  signal writePayloadToMem_buf_pointer :  std_logic_vector(35 downto 0);
  signal writePayloadToMem_packet_size_32 :  std_logic_vector(7 downto 0);
  signal writePayloadToMem_bad_packet_identifier :  std_logic_vector(0 downto 0);
  signal writePayloadToMem_last_keep :  std_logic_vector(7 downto 0);
  signal writePayloadToMem_in_args    : std_logic_vector(71 downto 0);
  signal writePayloadToMem_out_args   : std_logic_vector(16 downto 0);
  signal writePayloadToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writePayloadToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writePayloadToMem_start_req : std_logic;
  signal writePayloadToMem_start_ack : std_logic;
  signal writePayloadToMem_fin_req   : std_logic;
  signal writePayloadToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writePayloadToMem
  signal writePayloadToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writePayloadToMem_call_acks: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_acks: std_logic_vector(0 downto 0);
  signal writePayloadToMem_call_data: std_logic_vector(71 downto 0);
  signal writePayloadToMem_call_tag: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_data: std_logic_vector(16 downto 0);
  signal writePayloadToMem_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe AFB_NIC_REQUEST
  signal AFB_NIC_REQUEST_pipe_read_data: std_logic_vector(73 downto 0);
  signal AFB_NIC_REQUEST_pipe_read_req: std_logic_vector(0 downto 0);
  signal AFB_NIC_REQUEST_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe AFB_NIC_RESPONSE
  signal AFB_NIC_RESPONSE_pipe_write_data: std_logic_vector(32 downto 0);
  signal AFB_NIC_RESPONSE_pipe_write_req: std_logic_vector(0 downto 0);
  signal AFB_NIC_RESPONSE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe CONTROL_REGISTER
  signal CONTROL_REGISTER_pipe_write_data: std_logic_vector(31 downto 0);
  signal CONTROL_REGISTER_pipe_write_req: std_logic_vector(0 downto 0);
  signal CONTROL_REGISTER_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe CONTROL_REGISTER
  signal CONTROL_REGISTER: std_logic_vector(31 downto 0);
  -- aggregate signals for write to pipe FREE_Q
  signal FREE_Q_pipe_write_data: std_logic_vector(35 downto 0);
  signal FREE_Q_pipe_write_req: std_logic_vector(0 downto 0);
  signal FREE_Q_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe FREE_Q
  signal FREE_Q: std_logic_vector(35 downto 0);
  -- aggregate signals for write to pipe LAST_READ_TX_QUEUE_INDEX
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_data: std_logic_vector(11 downto 0);
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_req: std_logic_vector(1 downto 0);
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_ack: std_logic_vector(1 downto 0);
  -- signal decl. for read from internal signal pipe LAST_READ_TX_QUEUE_INDEX
  signal LAST_READ_TX_QUEUE_INDEX: std_logic_vector(5 downto 0);
  -- aggregate signals for write to pipe LAST_WRITTEN_RX_QUEUE_INDEX
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data: std_logic_vector(11 downto 0);
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req: std_logic_vector(1 downto 0);
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack: std_logic_vector(1 downto 0);
  -- signal decl. for read from internal signal pipe LAST_WRITTEN_RX_QUEUE_INDEX
  signal LAST_WRITTEN_RX_QUEUE_INDEX: std_logic_vector(5 downto 0);
  -- aggregate signals for read from pipe MEMORY_TO_NIC_RESPONSE
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_data: std_logic_vector(64 downto 0);
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_req: std_logic_vector(0 downto 0);
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_REQUEST_REGISTER_ACCESS_PIPE
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data: std_logic_vector(42 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe NIC_REQUEST_REGISTER_ACCESS_PIPE
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data: std_logic_vector(42 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req: std_logic_vector(0 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_RESPONSE_REGISTER_ACCESS_PIPE
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data: std_logic_vector(32 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe NIC_RESPONSE_REGISTER_ACCESS_PIPE
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data: std_logic_vector(32 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req: std_logic_vector(0 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_TO_MEMORY_REQUEST
  signal NIC_TO_MEMORY_REQUEST_pipe_write_data: std_logic_vector(109 downto 0);
  signal NIC_TO_MEMORY_REQUEST_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_TO_MEMORY_REQUEST_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NUMBER_OF_SERVERS
  signal NUMBER_OF_SERVERS_pipe_write_data: std_logic_vector(31 downto 0);
  signal NUMBER_OF_SERVERS_pipe_write_req: std_logic_vector(0 downto 0);
  signal NUMBER_OF_SERVERS_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe NUMBER_OF_SERVERS
  signal NUMBER_OF_SERVERS: std_logic_vector(31 downto 0);
  -- aggregate signals for read from pipe mac_to_nic_data
  signal mac_to_nic_data_pipe_read_data: std_logic_vector(72 downto 0);
  signal mac_to_nic_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal mac_to_nic_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_rx_to_header
  signal nic_rx_to_header_pipe_write_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_header_pipe_write_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_header_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe nic_rx_to_header
  signal nic_rx_to_header_pipe_read_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_header_pipe_read_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_header_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_rx_to_packet
  signal nic_rx_to_packet_pipe_write_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_packet_pipe_write_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_packet_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe nic_rx_to_packet
  signal nic_rx_to_packet_pipe_read_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_packet_pipe_read_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_packet_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_to_mac_transmit_pipe
  signal nic_to_mac_transmit_pipe_pipe_write_data: std_logic_vector(145 downto 0);
  signal nic_to_mac_transmit_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal nic_to_mac_transmit_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module AccessRegister
  AccessRegister_rwbar <= AccessRegister_in_args(42 downto 42);
  AccessRegister_bmask <= AccessRegister_in_args(41 downto 38);
  AccessRegister_register_index <= AccessRegister_in_args(37 downto 32);
  AccessRegister_wdata <= AccessRegister_in_args(31 downto 0);
  AccessRegister_out_args <= AccessRegister_rdata ;
  -- call arbiter for module AccessRegister
  AccessRegister_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 4,
      call_data_width => 43,
      return_data_width => 32,
      callee_tag_length => 3,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => AccessRegister_call_reqs,
      call_acks => AccessRegister_call_acks,
      return_reqs => AccessRegister_return_reqs,
      return_acks => AccessRegister_return_acks,
      call_data  => AccessRegister_call_data,
      call_tag  => AccessRegister_call_tag,
      return_tag  => AccessRegister_return_tag,
      call_mtag => AccessRegister_tag_in,
      return_mtag => AccessRegister_tag_out,
      return_data =>AccessRegister_return_data,
      call_mreq => AccessRegister_start_req,
      call_mack => AccessRegister_start_ack,
      return_mreq => AccessRegister_fin_req,
      return_mack => AccessRegister_fin_ack,
      call_mdata => AccessRegister_in_args,
      return_mdata => AccessRegister_out_args,
      clk => clk, 
      reset => reset --
    ); --
  AccessRegister_instance:AccessRegister-- 
    generic map(tag_length => 5)
    port map(-- 
      rwbar => AccessRegister_rwbar,
      bmask => AccessRegister_bmask,
      register_index => AccessRegister_register_index,
      wdata => AccessRegister_wdata,
      rdata => AccessRegister_rdata,
      start_req => AccessRegister_start_req,
      start_ack => AccessRegister_start_ack,
      fin_req => AccessRegister_fin_req,
      fin_ack => AccessRegister_fin_ack,
      clk => clk,
      reset => reset,
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data(32 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data(42 downto 0),
      tag_in => AccessRegister_tag_in,
      tag_out => AccessRegister_tag_out-- 
    ); -- 
  -- module NicRegisterAccessDaemon
  NicRegisterAccessDaemon_instance:NicRegisterAccessDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => NicRegisterAccessDaemon_start_req,
      start_ack => NicRegisterAccessDaemon_start_ack,
      fin_req => NicRegisterAccessDaemon_fin_req,
      fin_ack => NicRegisterAccessDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(11 downto 6),
      memory_space_0_lr_tag => memory_space_0_lr_tag(39 downto 20),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 32),
      memory_space_0_lc_tag => memory_space_0_lc_tag(5 downto 3),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data(42 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data(32 downto 0),
      UpdateRegister_call_reqs => UpdateRegister_call_reqs(1 downto 1),
      UpdateRegister_call_acks => UpdateRegister_call_acks(1 downto 1),
      UpdateRegister_call_data => UpdateRegister_call_data(147 downto 74),
      UpdateRegister_call_tag => UpdateRegister_call_tag(1 downto 1),
      UpdateRegister_return_reqs => UpdateRegister_return_reqs(1 downto 1),
      UpdateRegister_return_acks => UpdateRegister_return_acks(1 downto 1),
      UpdateRegister_return_data => UpdateRegister_return_data(63 downto 32),
      UpdateRegister_return_tag => UpdateRegister_return_tag(1 downto 1),
      tag_in => NicRegisterAccessDaemon_tag_in,
      tag_out => NicRegisterAccessDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  NicRegisterAccessDaemon_tag_in <= (others => '0');
  NicRegisterAccessDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => NicRegisterAccessDaemon_start_req, start_ack => NicRegisterAccessDaemon_start_ack,  fin_req => NicRegisterAccessDaemon_fin_req,  fin_ack => NicRegisterAccessDaemon_fin_ack);
  -- module ReceiveEngineDaemon
  ReceiveEngineDaemon_instance:ReceiveEngineDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => ReceiveEngineDaemon_start_req,
      start_ack => ReceiveEngineDaemon_start_ack,
      fin_req => ReceiveEngineDaemon_fin_req,
      fin_ack => ReceiveEngineDaemon_fin_ack,
      clk => clk,
      reset => reset,
      FREE_Q => FREE_Q,
      CONTROL_REGISTER => CONTROL_REGISTER,
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0 downto 0),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0 downto 0),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(5 downto 0),
      popFromQueue_call_reqs => popFromQueue_call_reqs(1 downto 1),
      popFromQueue_call_acks => popFromQueue_call_acks(1 downto 1),
      popFromQueue_call_data => popFromQueue_call_data(73 downto 37),
      popFromQueue_call_tag => popFromQueue_call_tag(1 downto 1),
      popFromQueue_return_reqs => popFromQueue_return_reqs(1 downto 1),
      popFromQueue_return_acks => popFromQueue_return_acks(1 downto 1),
      popFromQueue_return_data => popFromQueue_return_data(65 downto 33),
      popFromQueue_return_tag => popFromQueue_return_tag(1 downto 1),
      loadBuffer_call_reqs => loadBuffer_call_reqs(0 downto 0),
      loadBuffer_call_acks => loadBuffer_call_acks(0 downto 0),
      loadBuffer_call_data => loadBuffer_call_data(35 downto 0),
      loadBuffer_call_tag => loadBuffer_call_tag(0 downto 0),
      loadBuffer_return_reqs => loadBuffer_return_reqs(0 downto 0),
      loadBuffer_return_acks => loadBuffer_return_acks(0 downto 0),
      loadBuffer_return_data => loadBuffer_return_data(0 downto 0),
      loadBuffer_return_tag => loadBuffer_return_tag(0 downto 0),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(1 downto 1),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(1 downto 1),
      pushIntoQueue_call_data => pushIntoQueue_call_data(137 downto 69),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(1 downto 1),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(1 downto 1),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(1 downto 1),
      pushIntoQueue_return_data => pushIntoQueue_return_data(1 downto 1),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(1 downto 1),
      populateRxQueue_call_reqs => populateRxQueue_call_reqs(0 downto 0),
      populateRxQueue_call_acks => populateRxQueue_call_acks(0 downto 0),
      populateRxQueue_call_data => populateRxQueue_call_data(35 downto 0),
      populateRxQueue_call_tag => populateRxQueue_call_tag(0 downto 0),
      populateRxQueue_return_reqs => populateRxQueue_return_reqs(0 downto 0),
      populateRxQueue_return_acks => populateRxQueue_return_acks(0 downto 0),
      populateRxQueue_return_tag => populateRxQueue_return_tag(0 downto 0),
      tag_in => ReceiveEngineDaemon_tag_in,
      tag_out => ReceiveEngineDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  ReceiveEngineDaemon_tag_in <= (others => '0');
  ReceiveEngineDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ReceiveEngineDaemon_start_req, start_ack => ReceiveEngineDaemon_start_ack,  fin_req => ReceiveEngineDaemon_fin_req,  fin_ack => ReceiveEngineDaemon_fin_ack);
  -- module SoftwareRegisterAccessDaemon
  SoftwareRegisterAccessDaemon_instance:SoftwareRegisterAccessDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => SoftwareRegisterAccessDaemon_start_req,
      start_ack => SoftwareRegisterAccessDaemon_start_ack,
      fin_req => SoftwareRegisterAccessDaemon_fin_req,
      fin_ack => SoftwareRegisterAccessDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(5 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(19 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 0),
      AFB_NIC_REQUEST_pipe_read_req => AFB_NIC_REQUEST_pipe_read_req(0 downto 0),
      AFB_NIC_REQUEST_pipe_read_ack => AFB_NIC_REQUEST_pipe_read_ack(0 downto 0),
      AFB_NIC_REQUEST_pipe_read_data => AFB_NIC_REQUEST_pipe_read_data(73 downto 0),
      FREE_Q_pipe_write_req => FREE_Q_pipe_write_req(0 downto 0),
      FREE_Q_pipe_write_ack => FREE_Q_pipe_write_ack(0 downto 0),
      FREE_Q_pipe_write_data => FREE_Q_pipe_write_data(35 downto 0),
      AFB_NIC_RESPONSE_pipe_write_req => AFB_NIC_RESPONSE_pipe_write_req(0 downto 0),
      AFB_NIC_RESPONSE_pipe_write_ack => AFB_NIC_RESPONSE_pipe_write_ack(0 downto 0),
      AFB_NIC_RESPONSE_pipe_write_data => AFB_NIC_RESPONSE_pipe_write_data(32 downto 0),
      CONTROL_REGISTER_pipe_write_req => CONTROL_REGISTER_pipe_write_req(0 downto 0),
      CONTROL_REGISTER_pipe_write_ack => CONTROL_REGISTER_pipe_write_ack(0 downto 0),
      CONTROL_REGISTER_pipe_write_data => CONTROL_REGISTER_pipe_write_data(31 downto 0),
      NUMBER_OF_SERVERS_pipe_write_req => NUMBER_OF_SERVERS_pipe_write_req(0 downto 0),
      NUMBER_OF_SERVERS_pipe_write_ack => NUMBER_OF_SERVERS_pipe_write_ack(0 downto 0),
      NUMBER_OF_SERVERS_pipe_write_data => NUMBER_OF_SERVERS_pipe_write_data(31 downto 0),
      UpdateRegister_call_reqs => UpdateRegister_call_reqs(0 downto 0),
      UpdateRegister_call_acks => UpdateRegister_call_acks(0 downto 0),
      UpdateRegister_call_data => UpdateRegister_call_data(73 downto 0),
      UpdateRegister_call_tag => UpdateRegister_call_tag(0 downto 0),
      UpdateRegister_return_reqs => UpdateRegister_return_reqs(0 downto 0),
      UpdateRegister_return_acks => UpdateRegister_return_acks(0 downto 0),
      UpdateRegister_return_data => UpdateRegister_return_data(31 downto 0),
      UpdateRegister_return_tag => UpdateRegister_return_tag(0 downto 0),
      tag_in => SoftwareRegisterAccessDaemon_tag_in,
      tag_out => SoftwareRegisterAccessDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  SoftwareRegisterAccessDaemon_tag_in <= (others => '0');
  SoftwareRegisterAccessDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => SoftwareRegisterAccessDaemon_start_req, start_ack => SoftwareRegisterAccessDaemon_start_ack,  fin_req => SoftwareRegisterAccessDaemon_fin_req,  fin_ack => SoftwareRegisterAccessDaemon_fin_ack);
  -- module UpdateRegister
  UpdateRegister_bmask <= UpdateRegister_in_args(73 downto 70);
  UpdateRegister_rval <= UpdateRegister_in_args(69 downto 38);
  UpdateRegister_wdata <= UpdateRegister_in_args(37 downto 6);
  UpdateRegister_index <= UpdateRegister_in_args(5 downto 0);
  UpdateRegister_out_args <= UpdateRegister_wval ;
  -- call arbiter for module UpdateRegister
  UpdateRegister_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 74,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => UpdateRegister_call_reqs,
      call_acks => UpdateRegister_call_acks,
      return_reqs => UpdateRegister_return_reqs,
      return_acks => UpdateRegister_return_acks,
      call_data  => UpdateRegister_call_data,
      call_tag  => UpdateRegister_call_tag,
      return_tag  => UpdateRegister_return_tag,
      call_mtag => UpdateRegister_tag_in,
      return_mtag => UpdateRegister_tag_out,
      return_data =>UpdateRegister_return_data,
      call_mreq => UpdateRegister_start_req,
      call_mack => UpdateRegister_start_ack,
      return_mreq => UpdateRegister_fin_req,
      return_mack => UpdateRegister_fin_ack,
      call_mdata => UpdateRegister_in_args,
      return_mdata => UpdateRegister_out_args,
      clk => clk, 
      reset => reset --
    ); --
  UpdateRegister_instance:UpdateRegister-- 
    generic map(tag_length => 3)
    port map(-- 
      bmask => UpdateRegister_bmask,
      rval => UpdateRegister_rval,
      wdata => UpdateRegister_wdata,
      index => UpdateRegister_index,
      wval => UpdateRegister_wval,
      start_req => UpdateRegister_start_req,
      start_ack => UpdateRegister_start_ack,
      fin_req => UpdateRegister_fin_req,
      fin_ack => UpdateRegister_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(5 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(31 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(19 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(2 downto 0),
      tag_in => UpdateRegister_tag_in,
      tag_out => UpdateRegister_tag_out-- 
    ); -- 
  -- module accessMemory
  accessMemory_lock <= accessMemory_in_args(109 downto 109);
  accessMemory_rwbar <= accessMemory_in_args(108 downto 108);
  accessMemory_bmask <= accessMemory_in_args(107 downto 100);
  accessMemory_addr <= accessMemory_in_args(99 downto 64);
  accessMemory_wdata <= accessMemory_in_args(63 downto 0);
  accessMemory_out_args <= accessMemory_rdata ;
  -- call arbiter for module accessMemory
  accessMemory_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 11,
      call_data_width => 110,
      return_data_width => 64,
      callee_tag_length => 4,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => accessMemory_call_reqs,
      call_acks => accessMemory_call_acks,
      return_reqs => accessMemory_return_reqs,
      return_acks => accessMemory_return_acks,
      call_data  => accessMemory_call_data,
      call_tag  => accessMemory_call_tag,
      return_tag  => accessMemory_return_tag,
      call_mtag => accessMemory_tag_in,
      return_mtag => accessMemory_tag_out,
      return_data =>accessMemory_return_data,
      call_mreq => accessMemory_start_req,
      call_mack => accessMemory_start_ack,
      return_mreq => accessMemory_fin_req,
      return_mack => accessMemory_fin_ack,
      call_mdata => accessMemory_in_args,
      return_mdata => accessMemory_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMemory_instance:accessMemory-- 
    generic map(tag_length => 6)
    port map(-- 
      lock => accessMemory_lock,
      rwbar => accessMemory_rwbar,
      bmask => accessMemory_bmask,
      addr => accessMemory_addr,
      wdata => accessMemory_wdata,
      rdata => accessMemory_rdata,
      start_req => accessMemory_start_req,
      start_ack => accessMemory_start_ack,
      fin_req => accessMemory_fin_req,
      fin_ack => accessMemory_fin_ack,
      clk => clk,
      reset => reset,
      MEMORY_TO_NIC_RESPONSE_pipe_read_req => MEMORY_TO_NIC_RESPONSE_pipe_read_req(0 downto 0),
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack(0 downto 0),
      MEMORY_TO_NIC_RESPONSE_pipe_read_data => MEMORY_TO_NIC_RESPONSE_pipe_read_data(64 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_req => NIC_TO_MEMORY_REQUEST_pipe_write_req(0 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_ack => NIC_TO_MEMORY_REQUEST_pipe_write_ack(0 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_data => NIC_TO_MEMORY_REQUEST_pipe_write_data(109 downto 0),
      tag_in => accessMemory_tag_in,
      tag_out => accessMemory_tag_out-- 
    ); -- 
  -- module acquireMutex
  acquireMutex_q_base_address <= acquireMutex_in_args(35 downto 0);
  acquireMutex_out_args <= acquireMutex_m_ok ;
  -- call arbiter for module acquireMutex
  acquireMutex_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 36,
      return_data_width => 1,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => acquireMutex_call_reqs,
      call_acks => acquireMutex_call_acks,
      return_reqs => acquireMutex_return_reqs,
      return_acks => acquireMutex_return_acks,
      call_data  => acquireMutex_call_data,
      call_tag  => acquireMutex_call_tag,
      return_tag  => acquireMutex_return_tag,
      call_mtag => acquireMutex_tag_in,
      return_mtag => acquireMutex_tag_out,
      return_data =>acquireMutex_return_data,
      call_mreq => acquireMutex_start_req,
      call_mack => acquireMutex_start_ack,
      return_mreq => acquireMutex_fin_req,
      return_mack => acquireMutex_fin_ack,
      call_mdata => acquireMutex_in_args,
      return_mdata => acquireMutex_out_args,
      clk => clk, 
      reset => reset --
    ); --
  acquireMutex_instance:acquireMutex-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => acquireMutex_q_base_address,
      m_ok => acquireMutex_m_ok,
      start_req => acquireMutex_start_req,
      start_ack => acquireMutex_start_ack,
      fin_req => acquireMutex_fin_req,
      fin_ack => acquireMutex_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(6 downto 6),
      accessMemory_call_acks => accessMemory_call_acks(6 downto 6),
      accessMemory_call_data => accessMemory_call_data(769 downto 660),
      accessMemory_call_tag => accessMemory_call_tag(13 downto 12),
      accessMemory_return_reqs => accessMemory_return_reqs(6 downto 6),
      accessMemory_return_acks => accessMemory_return_acks(6 downto 6),
      accessMemory_return_data => accessMemory_return_data(447 downto 384),
      accessMemory_return_tag => accessMemory_return_tag(13 downto 12),
      tag_in => acquireMutex_tag_in,
      tag_out => acquireMutex_tag_out-- 
    ); -- 
  -- module getQueueElement
  getQueueElement_q_base_address <= getQueueElement_in_args(67 downto 32);
  getQueueElement_read_pointer <= getQueueElement_in_args(31 downto 0);
  getQueueElement_out_args <= getQueueElement_q_r_data ;
  -- call arbiter for module getQueueElement
  getQueueElement_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 68,
      return_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueueElement_call_reqs,
      call_acks => getQueueElement_call_acks,
      return_reqs => getQueueElement_return_reqs,
      return_acks => getQueueElement_return_acks,
      call_data  => getQueueElement_call_data,
      call_tag  => getQueueElement_call_tag,
      return_tag  => getQueueElement_return_tag,
      call_mtag => getQueueElement_tag_in,
      return_mtag => getQueueElement_tag_out,
      return_data =>getQueueElement_return_data,
      call_mreq => getQueueElement_start_req,
      call_mack => getQueueElement_start_ack,
      return_mreq => getQueueElement_fin_req,
      return_mack => getQueueElement_fin_ack,
      call_mdata => getQueueElement_in_args,
      return_mdata => getQueueElement_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueueElement_instance:getQueueElement-- 
    generic map(tag_length => 2)
    port map(-- 
      q_base_address => getQueueElement_q_base_address,
      read_pointer => getQueueElement_read_pointer,
      q_r_data => getQueueElement_q_r_data,
      start_req => getQueueElement_start_req,
      start_ack => getQueueElement_start_ack,
      fin_req => getQueueElement_fin_req,
      fin_ack => getQueueElement_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(7 downto 7),
      accessMemory_call_acks => accessMemory_call_acks(7 downto 7),
      accessMemory_call_data => accessMemory_call_data(879 downto 770),
      accessMemory_call_tag => accessMemory_call_tag(15 downto 14),
      accessMemory_return_reqs => accessMemory_return_reqs(7 downto 7),
      accessMemory_return_acks => accessMemory_return_acks(7 downto 7),
      accessMemory_return_data => accessMemory_return_data(511 downto 448),
      accessMemory_return_tag => accessMemory_return_tag(15 downto 14),
      tag_in => getQueueElement_tag_in,
      tag_out => getQueueElement_tag_out-- 
    ); -- 
  -- module getQueuePointers
  getQueuePointers_q_base_address <= getQueuePointers_in_args(35 downto 0);
  getQueuePointers_out_args <= getQueuePointers_wp & getQueuePointers_rp ;
  -- call arbiter for module getQueuePointers
  getQueuePointers_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 36,
      return_data_width => 64,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueuePointers_call_reqs,
      call_acks => getQueuePointers_call_acks,
      return_reqs => getQueuePointers_return_reqs,
      return_acks => getQueuePointers_return_acks,
      call_data  => getQueuePointers_call_data,
      call_tag  => getQueuePointers_call_tag,
      return_tag  => getQueuePointers_return_tag,
      call_mtag => getQueuePointers_tag_in,
      return_mtag => getQueuePointers_tag_out,
      return_data =>getQueuePointers_return_data,
      call_mreq => getQueuePointers_start_req,
      call_mack => getQueuePointers_start_ack,
      return_mreq => getQueuePointers_fin_req,
      return_mack => getQueuePointers_fin_ack,
      call_mdata => getQueuePointers_in_args,
      return_mdata => getQueuePointers_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueuePointers_instance:getQueuePointers-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => getQueuePointers_q_base_address,
      wp => getQueuePointers_wp,
      rp => getQueuePointers_rp,
      start_req => getQueuePointers_start_req,
      start_ack => getQueuePointers_start_ack,
      fin_req => getQueuePointers_fin_req,
      fin_ack => getQueuePointers_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(8 downto 8),
      accessMemory_call_acks => accessMemory_call_acks(8 downto 8),
      accessMemory_call_data => accessMemory_call_data(989 downto 880),
      accessMemory_call_tag => accessMemory_call_tag(17 downto 16),
      accessMemory_return_reqs => accessMemory_return_reqs(8 downto 8),
      accessMemory_return_acks => accessMemory_return_acks(8 downto 8),
      accessMemory_return_data => accessMemory_return_data(575 downto 512),
      accessMemory_return_tag => accessMemory_return_tag(17 downto 16),
      tag_in => getQueuePointers_tag_in,
      tag_out => getQueuePointers_tag_out-- 
    ); -- 
  -- module getTxPacketPointerFromServer
  getTxPacketPointerFromServer_queue_index <= getTxPacketPointerFromServer_in_args(5 downto 0);
  getTxPacketPointerFromServer_out_args <= getTxPacketPointerFromServer_pkt_pointer & getTxPacketPointerFromServer_status ;
  -- call arbiter for module getTxPacketPointerFromServer
  getTxPacketPointerFromServer_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 6,
      return_data_width => 33,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getTxPacketPointerFromServer_call_reqs,
      call_acks => getTxPacketPointerFromServer_call_acks,
      return_reqs => getTxPacketPointerFromServer_return_reqs,
      return_acks => getTxPacketPointerFromServer_return_acks,
      call_data  => getTxPacketPointerFromServer_call_data,
      call_tag  => getTxPacketPointerFromServer_call_tag,
      return_tag  => getTxPacketPointerFromServer_return_tag,
      call_mtag => getTxPacketPointerFromServer_tag_in,
      return_mtag => getTxPacketPointerFromServer_tag_out,
      return_data =>getTxPacketPointerFromServer_return_data,
      call_mreq => getTxPacketPointerFromServer_start_req,
      call_mack => getTxPacketPointerFromServer_start_ack,
      return_mreq => getTxPacketPointerFromServer_fin_req,
      return_mack => getTxPacketPointerFromServer_fin_ack,
      call_mdata => getTxPacketPointerFromServer_in_args,
      return_mdata => getTxPacketPointerFromServer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getTxPacketPointerFromServer_instance:getTxPacketPointerFromServer-- 
    generic map(tag_length => 2)
    port map(-- 
      queue_index => getTxPacketPointerFromServer_queue_index,
      pkt_pointer => getTxPacketPointerFromServer_pkt_pointer,
      status => getTxPacketPointerFromServer_status,
      start_req => getTxPacketPointerFromServer_start_req,
      start_ack => getTxPacketPointerFromServer_start_ack,
      fin_req => getTxPacketPointerFromServer_fin_req,
      fin_ack => getTxPacketPointerFromServer_fin_ack,
      clk => clk,
      reset => reset,
      AccessRegister_call_reqs => AccessRegister_call_reqs(2 downto 2),
      AccessRegister_call_acks => AccessRegister_call_acks(2 downto 2),
      AccessRegister_call_data => AccessRegister_call_data(128 downto 86),
      AccessRegister_call_tag => AccessRegister_call_tag(5 downto 4),
      AccessRegister_return_reqs => AccessRegister_return_reqs(2 downto 2),
      AccessRegister_return_acks => AccessRegister_return_acks(2 downto 2),
      AccessRegister_return_data => AccessRegister_return_data(95 downto 64),
      AccessRegister_return_tag => AccessRegister_return_tag(5 downto 4),
      popFromQueue_call_reqs => popFromQueue_call_reqs(0 downto 0),
      popFromQueue_call_acks => popFromQueue_call_acks(0 downto 0),
      popFromQueue_call_data => popFromQueue_call_data(36 downto 0),
      popFromQueue_call_tag => popFromQueue_call_tag(0 downto 0),
      popFromQueue_return_reqs => popFromQueue_return_reqs(0 downto 0),
      popFromQueue_return_acks => popFromQueue_return_acks(0 downto 0),
      popFromQueue_return_data => popFromQueue_return_data(32 downto 0),
      popFromQueue_return_tag => popFromQueue_return_tag(0 downto 0),
      tag_in => getTxPacketPointerFromServer_tag_in,
      tag_out => getTxPacketPointerFromServer_tag_out-- 
    ); -- 
  -- module loadBuffer
  loadBuffer_rx_buffer_pointer <= loadBuffer_in_args(35 downto 0);
  loadBuffer_out_args <= loadBuffer_bad_packet_identifier ;
  -- call arbiter for module loadBuffer
  loadBuffer_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 36,
      return_data_width => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadBuffer_call_reqs,
      call_acks => loadBuffer_call_acks,
      return_reqs => loadBuffer_return_reqs,
      return_acks => loadBuffer_return_acks,
      call_data  => loadBuffer_call_data,
      call_tag  => loadBuffer_call_tag,
      return_tag  => loadBuffer_return_tag,
      call_mtag => loadBuffer_tag_in,
      return_mtag => loadBuffer_tag_out,
      return_data =>loadBuffer_return_data,
      call_mreq => loadBuffer_start_req,
      call_mack => loadBuffer_start_ack,
      return_mreq => loadBuffer_fin_req,
      return_mack => loadBuffer_fin_ack,
      call_mdata => loadBuffer_in_args,
      return_mdata => loadBuffer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  loadBuffer_instance:loadBuffer-- 
    generic map(tag_length => 2)
    port map(-- 
      rx_buffer_pointer => loadBuffer_rx_buffer_pointer,
      bad_packet_identifier => loadBuffer_bad_packet_identifier,
      start_req => loadBuffer_start_req,
      start_ack => loadBuffer_start_ack,
      fin_req => loadBuffer_fin_req,
      fin_ack => loadBuffer_fin_ack,
      clk => clk,
      reset => reset,
      writeEthernetHeaderToMem_call_reqs => writeEthernetHeaderToMem_call_reqs(0 downto 0),
      writeEthernetHeaderToMem_call_acks => writeEthernetHeaderToMem_call_acks(0 downto 0),
      writeEthernetHeaderToMem_call_data => writeEthernetHeaderToMem_call_data(35 downto 0),
      writeEthernetHeaderToMem_call_tag => writeEthernetHeaderToMem_call_tag(0 downto 0),
      writeEthernetHeaderToMem_return_reqs => writeEthernetHeaderToMem_return_reqs(0 downto 0),
      writeEthernetHeaderToMem_return_acks => writeEthernetHeaderToMem_return_acks(0 downto 0),
      writeEthernetHeaderToMem_return_data => writeEthernetHeaderToMem_return_data(35 downto 0),
      writeEthernetHeaderToMem_return_tag => writeEthernetHeaderToMem_return_tag(0 downto 0),
      writePayloadToMem_call_reqs => writePayloadToMem_call_reqs(0 downto 0),
      writePayloadToMem_call_acks => writePayloadToMem_call_acks(0 downto 0),
      writePayloadToMem_call_data => writePayloadToMem_call_data(71 downto 0),
      writePayloadToMem_call_tag => writePayloadToMem_call_tag(0 downto 0),
      writePayloadToMem_return_reqs => writePayloadToMem_return_reqs(0 downto 0),
      writePayloadToMem_return_acks => writePayloadToMem_return_acks(0 downto 0),
      writePayloadToMem_return_data => writePayloadToMem_return_data(16 downto 0),
      writePayloadToMem_return_tag => writePayloadToMem_return_tag(0 downto 0),
      writeControlInformationToMem_call_reqs => writeControlInformationToMem_call_reqs(0 downto 0),
      writeControlInformationToMem_call_acks => writeControlInformationToMem_call_acks(0 downto 0),
      writeControlInformationToMem_call_data => writeControlInformationToMem_call_data(51 downto 0),
      writeControlInformationToMem_call_tag => writeControlInformationToMem_call_tag(0 downto 0),
      writeControlInformationToMem_return_reqs => writeControlInformationToMem_return_reqs(0 downto 0),
      writeControlInformationToMem_return_acks => writeControlInformationToMem_return_acks(0 downto 0),
      writeControlInformationToMem_return_tag => writeControlInformationToMem_return_tag(0 downto 0),
      tag_in => loadBuffer_tag_in,
      tag_out => loadBuffer_tag_out-- 
    ); -- 
  -- module nicRxFromMacDaemon
  nicRxFromMacDaemon_instance:nicRxFromMacDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => nicRxFromMacDaemon_start_req,
      start_ack => nicRxFromMacDaemon_start_ack,
      fin_req => nicRxFromMacDaemon_fin_req,
      fin_ack => nicRxFromMacDaemon_fin_ack,
      clk => clk,
      reset => reset,
      CONTROL_REGISTER => CONTROL_REGISTER,
      mac_to_nic_data_pipe_read_req => mac_to_nic_data_pipe_read_req(0 downto 0),
      mac_to_nic_data_pipe_read_ack => mac_to_nic_data_pipe_read_ack(0 downto 0),
      mac_to_nic_data_pipe_read_data => mac_to_nic_data_pipe_read_data(72 downto 0),
      nic_rx_to_packet_pipe_write_req => nic_rx_to_packet_pipe_write_req(0 downto 0),
      nic_rx_to_packet_pipe_write_ack => nic_rx_to_packet_pipe_write_ack(0 downto 0),
      nic_rx_to_packet_pipe_write_data => nic_rx_to_packet_pipe_write_data(72 downto 0),
      nic_rx_to_header_pipe_write_req => nic_rx_to_header_pipe_write_req(0 downto 0),
      nic_rx_to_header_pipe_write_ack => nic_rx_to_header_pipe_write_ack(0 downto 0),
      nic_rx_to_header_pipe_write_data => nic_rx_to_header_pipe_write_data(72 downto 0),
      AccessRegister_call_reqs => AccessRegister_call_reqs(1 downto 1),
      AccessRegister_call_acks => AccessRegister_call_acks(1 downto 1),
      AccessRegister_call_data => AccessRegister_call_data(85 downto 43),
      AccessRegister_call_tag => AccessRegister_call_tag(3 downto 2),
      AccessRegister_return_reqs => AccessRegister_return_reqs(1 downto 1),
      AccessRegister_return_acks => AccessRegister_return_acks(1 downto 1),
      AccessRegister_return_data => AccessRegister_return_data(63 downto 32),
      AccessRegister_return_tag => AccessRegister_return_tag(3 downto 2),
      tag_in => nicRxFromMacDaemon_tag_in,
      tag_out => nicRxFromMacDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  nicRxFromMacDaemon_tag_in <= (others => '0');
  nicRxFromMacDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => nicRxFromMacDaemon_start_req, start_ack => nicRxFromMacDaemon_start_ack,  fin_req => nicRxFromMacDaemon_fin_req,  fin_ack => nicRxFromMacDaemon_fin_ack);
  -- module popFromQueue
  popFromQueue_lock <= popFromQueue_in_args(36 downto 36);
  popFromQueue_q_base_address <= popFromQueue_in_args(35 downto 0);
  popFromQueue_out_args <= popFromQueue_q_r_data & popFromQueue_status ;
  -- call arbiter for module popFromQueue
  popFromQueue_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 37,
      return_data_width => 33,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => popFromQueue_call_reqs,
      call_acks => popFromQueue_call_acks,
      return_reqs => popFromQueue_return_reqs,
      return_acks => popFromQueue_return_acks,
      call_data  => popFromQueue_call_data,
      call_tag  => popFromQueue_call_tag,
      return_tag  => popFromQueue_return_tag,
      call_mtag => popFromQueue_tag_in,
      return_mtag => popFromQueue_tag_out,
      return_data =>popFromQueue_return_data,
      call_mreq => popFromQueue_start_req,
      call_mack => popFromQueue_start_ack,
      return_mreq => popFromQueue_fin_req,
      return_mack => popFromQueue_fin_ack,
      call_mdata => popFromQueue_in_args,
      return_mdata => popFromQueue_out_args,
      clk => clk, 
      reset => reset --
    ); --
  popFromQueue_instance:popFromQueue-- 
    generic map(tag_length => 3)
    port map(-- 
      lock => popFromQueue_lock,
      q_base_address => popFromQueue_q_base_address,
      q_r_data => popFromQueue_q_r_data,
      status => popFromQueue_status,
      start_req => popFromQueue_start_req,
      start_ack => popFromQueue_start_ack,
      fin_req => popFromQueue_fin_req,
      fin_ack => popFromQueue_fin_ack,
      clk => clk,
      reset => reset,
      acquireMutex_call_reqs => acquireMutex_call_reqs(1 downto 1),
      acquireMutex_call_acks => acquireMutex_call_acks(1 downto 1),
      acquireMutex_call_data => acquireMutex_call_data(71 downto 36),
      acquireMutex_call_tag => acquireMutex_call_tag(1 downto 1),
      acquireMutex_return_reqs => acquireMutex_return_reqs(1 downto 1),
      acquireMutex_return_acks => acquireMutex_return_acks(1 downto 1),
      acquireMutex_return_data => acquireMutex_return_data(1 downto 1),
      acquireMutex_return_tag => acquireMutex_return_tag(1 downto 1),
      getQueuePointers_call_reqs => getQueuePointers_call_reqs(1 downto 1),
      getQueuePointers_call_acks => getQueuePointers_call_acks(1 downto 1),
      getQueuePointers_call_data => getQueuePointers_call_data(71 downto 36),
      getQueuePointers_call_tag => getQueuePointers_call_tag(1 downto 1),
      getQueuePointers_return_reqs => getQueuePointers_return_reqs(1 downto 1),
      getQueuePointers_return_acks => getQueuePointers_return_acks(1 downto 1),
      getQueuePointers_return_data => getQueuePointers_return_data(127 downto 64),
      getQueuePointers_return_tag => getQueuePointers_return_tag(1 downto 1),
      getQueueElement_call_reqs => getQueueElement_call_reqs(0 downto 0),
      getQueueElement_call_acks => getQueueElement_call_acks(0 downto 0),
      getQueueElement_call_data => getQueueElement_call_data(67 downto 0),
      getQueueElement_call_tag => getQueueElement_call_tag(0 downto 0),
      getQueueElement_return_reqs => getQueueElement_return_reqs(0 downto 0),
      getQueueElement_return_acks => getQueueElement_return_acks(0 downto 0),
      getQueueElement_return_data => getQueueElement_return_data(31 downto 0),
      getQueueElement_return_tag => getQueueElement_return_tag(0 downto 0),
      setQueuePointers_call_reqs => setQueuePointers_call_reqs(1 downto 1),
      setQueuePointers_call_acks => setQueuePointers_call_acks(1 downto 1),
      setQueuePointers_call_data => setQueuePointers_call_data(199 downto 100),
      setQueuePointers_call_tag => setQueuePointers_call_tag(1 downto 1),
      setQueuePointers_return_reqs => setQueuePointers_return_reqs(1 downto 1),
      setQueuePointers_return_acks => setQueuePointers_return_acks(1 downto 1),
      setQueuePointers_return_tag => setQueuePointers_return_tag(1 downto 1),
      releaseMutex_call_reqs => releaseMutex_call_reqs(1 downto 1),
      releaseMutex_call_acks => releaseMutex_call_acks(1 downto 1),
      releaseMutex_call_data => releaseMutex_call_data(71 downto 36),
      releaseMutex_call_tag => releaseMutex_call_tag(1 downto 1),
      releaseMutex_return_reqs => releaseMutex_return_reqs(1 downto 1),
      releaseMutex_return_acks => releaseMutex_return_acks(1 downto 1),
      releaseMutex_return_tag => releaseMutex_return_tag(1 downto 1),
      tag_in => popFromQueue_tag_in,
      tag_out => popFromQueue_tag_out-- 
    ); -- 
  -- module populateRxQueue
  populateRxQueue_rx_buffer_pointer <= populateRxQueue_in_args(35 downto 0);
  -- call arbiter for module populateRxQueue
  populateRxQueue_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 36,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => populateRxQueue_call_reqs,
      call_acks => populateRxQueue_call_acks,
      return_reqs => populateRxQueue_return_reqs,
      return_acks => populateRxQueue_return_acks,
      call_data  => populateRxQueue_call_data,
      call_tag  => populateRxQueue_call_tag,
      return_tag  => populateRxQueue_return_tag,
      call_mtag => populateRxQueue_tag_in,
      return_mtag => populateRxQueue_tag_out,
      call_mreq => populateRxQueue_start_req,
      call_mack => populateRxQueue_start_ack,
      return_mreq => populateRxQueue_fin_req,
      return_mack => populateRxQueue_fin_ack,
      call_mdata => populateRxQueue_in_args,
      clk => clk, 
      reset => reset --
    ); --
  populateRxQueue_instance:populateRxQueue-- 
    generic map(tag_length => 2)
    port map(-- 
      rx_buffer_pointer => populateRxQueue_rx_buffer_pointer,
      start_req => populateRxQueue_start_req,
      start_ack => populateRxQueue_start_ack,
      fin_req => populateRxQueue_fin_req,
      fin_ack => populateRxQueue_fin_ack,
      clk => clk,
      reset => reset,
      LAST_WRITTEN_RX_QUEUE_INDEX => LAST_WRITTEN_RX_QUEUE_INDEX,
      NUMBER_OF_SERVERS => NUMBER_OF_SERVERS,
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(1 downto 1),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(1 downto 1),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(11 downto 6),
      AccessRegister_call_reqs => AccessRegister_call_reqs(3 downto 3),
      AccessRegister_call_acks => AccessRegister_call_acks(3 downto 3),
      AccessRegister_call_data => AccessRegister_call_data(171 downto 129),
      AccessRegister_call_tag => AccessRegister_call_tag(7 downto 6),
      AccessRegister_return_reqs => AccessRegister_return_reqs(3 downto 3),
      AccessRegister_return_acks => AccessRegister_return_acks(3 downto 3),
      AccessRegister_return_data => AccessRegister_return_data(127 downto 96),
      AccessRegister_return_tag => AccessRegister_return_tag(7 downto 6),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(2 downto 2),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(2 downto 2),
      pushIntoQueue_call_data => pushIntoQueue_call_data(206 downto 138),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(2 downto 2),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(2 downto 2),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(2 downto 2),
      pushIntoQueue_return_data => pushIntoQueue_return_data(2 downto 2),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(2 downto 2),
      tag_in => populateRxQueue_tag_in,
      tag_out => populateRxQueue_tag_out-- 
    ); -- 
  -- module pushIntoQueue
  pushIntoQueue_lock <= pushIntoQueue_in_args(68 downto 68);
  pushIntoQueue_q_base_address <= pushIntoQueue_in_args(67 downto 32);
  pushIntoQueue_q_w_data <= pushIntoQueue_in_args(31 downto 0);
  pushIntoQueue_out_args <= pushIntoQueue_status ;
  -- call arbiter for module pushIntoQueue
  pushIntoQueue_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 3,
      call_data_width => 69,
      return_data_width => 1,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => pushIntoQueue_call_reqs,
      call_acks => pushIntoQueue_call_acks,
      return_reqs => pushIntoQueue_return_reqs,
      return_acks => pushIntoQueue_return_acks,
      call_data  => pushIntoQueue_call_data,
      call_tag  => pushIntoQueue_call_tag,
      return_tag  => pushIntoQueue_return_tag,
      call_mtag => pushIntoQueue_tag_in,
      return_mtag => pushIntoQueue_tag_out,
      return_data =>pushIntoQueue_return_data,
      call_mreq => pushIntoQueue_start_req,
      call_mack => pushIntoQueue_start_ack,
      return_mreq => pushIntoQueue_fin_req,
      return_mack => pushIntoQueue_fin_ack,
      call_mdata => pushIntoQueue_in_args,
      return_mdata => pushIntoQueue_out_args,
      clk => clk, 
      reset => reset --
    ); --
  pushIntoQueue_instance:pushIntoQueue-- 
    generic map(tag_length => 3)
    port map(-- 
      lock => pushIntoQueue_lock,
      q_base_address => pushIntoQueue_q_base_address,
      q_w_data => pushIntoQueue_q_w_data,
      status => pushIntoQueue_status,
      start_req => pushIntoQueue_start_req,
      start_ack => pushIntoQueue_start_ack,
      fin_req => pushIntoQueue_fin_req,
      fin_ack => pushIntoQueue_fin_ack,
      clk => clk,
      reset => reset,
      acquireMutex_call_reqs => acquireMutex_call_reqs(0 downto 0),
      acquireMutex_call_acks => acquireMutex_call_acks(0 downto 0),
      acquireMutex_call_data => acquireMutex_call_data(35 downto 0),
      acquireMutex_call_tag => acquireMutex_call_tag(0 downto 0),
      acquireMutex_return_reqs => acquireMutex_return_reqs(0 downto 0),
      acquireMutex_return_acks => acquireMutex_return_acks(0 downto 0),
      acquireMutex_return_data => acquireMutex_return_data(0 downto 0),
      acquireMutex_return_tag => acquireMutex_return_tag(0 downto 0),
      getQueuePointers_call_reqs => getQueuePointers_call_reqs(0 downto 0),
      getQueuePointers_call_acks => getQueuePointers_call_acks(0 downto 0),
      getQueuePointers_call_data => getQueuePointers_call_data(35 downto 0),
      getQueuePointers_call_tag => getQueuePointers_call_tag(0 downto 0),
      getQueuePointers_return_reqs => getQueuePointers_return_reqs(0 downto 0),
      getQueuePointers_return_acks => getQueuePointers_return_acks(0 downto 0),
      getQueuePointers_return_data => getQueuePointers_return_data(63 downto 0),
      getQueuePointers_return_tag => getQueuePointers_return_tag(0 downto 0),
      setQueuePointers_call_reqs => setQueuePointers_call_reqs(0 downto 0),
      setQueuePointers_call_acks => setQueuePointers_call_acks(0 downto 0),
      setQueuePointers_call_data => setQueuePointers_call_data(99 downto 0),
      setQueuePointers_call_tag => setQueuePointers_call_tag(0 downto 0),
      setQueuePointers_return_reqs => setQueuePointers_return_reqs(0 downto 0),
      setQueuePointers_return_acks => setQueuePointers_return_acks(0 downto 0),
      setQueuePointers_return_tag => setQueuePointers_return_tag(0 downto 0),
      releaseMutex_call_reqs => releaseMutex_call_reqs(0 downto 0),
      releaseMutex_call_acks => releaseMutex_call_acks(0 downto 0),
      releaseMutex_call_data => releaseMutex_call_data(35 downto 0),
      releaseMutex_call_tag => releaseMutex_call_tag(0 downto 0),
      releaseMutex_return_reqs => releaseMutex_return_reqs(0 downto 0),
      releaseMutex_return_acks => releaseMutex_return_acks(0 downto 0),
      releaseMutex_return_tag => releaseMutex_return_tag(0 downto 0),
      setQueueElement_call_reqs => setQueueElement_call_reqs(0 downto 0),
      setQueueElement_call_acks => setQueueElement_call_acks(0 downto 0),
      setQueueElement_call_data => setQueueElement_call_data(99 downto 0),
      setQueueElement_call_tag => setQueueElement_call_tag(0 downto 0),
      setQueueElement_return_reqs => setQueueElement_return_reqs(0 downto 0),
      setQueueElement_return_acks => setQueueElement_return_acks(0 downto 0),
      setQueueElement_return_tag => setQueueElement_return_tag(0 downto 0),
      tag_in => pushIntoQueue_tag_in,
      tag_out => pushIntoQueue_tag_out-- 
    ); -- 
  -- module releaseMutex
  releaseMutex_q_base_address <= releaseMutex_in_args(35 downto 0);
  -- call arbiter for module releaseMutex
  releaseMutex_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 2,
      call_data_width => 36,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => releaseMutex_call_reqs,
      call_acks => releaseMutex_call_acks,
      return_reqs => releaseMutex_return_reqs,
      return_acks => releaseMutex_return_acks,
      call_data  => releaseMutex_call_data,
      call_tag  => releaseMutex_call_tag,
      return_tag  => releaseMutex_return_tag,
      call_mtag => releaseMutex_tag_in,
      return_mtag => releaseMutex_tag_out,
      call_mreq => releaseMutex_start_req,
      call_mack => releaseMutex_start_ack,
      return_mreq => releaseMutex_fin_req,
      return_mack => releaseMutex_fin_ack,
      call_mdata => releaseMutex_in_args,
      clk => clk, 
      reset => reset --
    ); --
  releaseMutex_instance:releaseMutex-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => releaseMutex_q_base_address,
      start_req => releaseMutex_start_req,
      start_ack => releaseMutex_start_ack,
      fin_req => releaseMutex_fin_req,
      fin_ack => releaseMutex_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(9 downto 9),
      accessMemory_call_acks => accessMemory_call_acks(9 downto 9),
      accessMemory_call_data => accessMemory_call_data(1099 downto 990),
      accessMemory_call_tag => accessMemory_call_tag(19 downto 18),
      accessMemory_return_reqs => accessMemory_return_reqs(9 downto 9),
      accessMemory_return_acks => accessMemory_return_acks(9 downto 9),
      accessMemory_return_data => accessMemory_return_data(639 downto 576),
      accessMemory_return_tag => accessMemory_return_tag(19 downto 18),
      tag_in => releaseMutex_tag_in,
      tag_out => releaseMutex_tag_out-- 
    ); -- 
  -- module setQueueElement
  setQueueElement_q_base_address <= setQueueElement_in_args(99 downto 64);
  setQueueElement_write_pointer <= setQueueElement_in_args(63 downto 32);
  setQueueElement_q_w_data <= setQueueElement_in_args(31 downto 0);
  -- call arbiter for module setQueueElement
  setQueueElement_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 100,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => setQueueElement_call_reqs,
      call_acks => setQueueElement_call_acks,
      return_reqs => setQueueElement_return_reqs,
      return_acks => setQueueElement_return_acks,
      call_data  => setQueueElement_call_data,
      call_tag  => setQueueElement_call_tag,
      return_tag  => setQueueElement_return_tag,
      call_mtag => setQueueElement_tag_in,
      return_mtag => setQueueElement_tag_out,
      call_mreq => setQueueElement_start_req,
      call_mack => setQueueElement_start_ack,
      return_mreq => setQueueElement_fin_req,
      return_mack => setQueueElement_fin_ack,
      call_mdata => setQueueElement_in_args,
      clk => clk, 
      reset => reset --
    ); --
  setQueueElement_instance:setQueueElement-- 
    generic map(tag_length => 2)
    port map(-- 
      q_base_address => setQueueElement_q_base_address,
      write_pointer => setQueueElement_write_pointer,
      q_w_data => setQueueElement_q_w_data,
      start_req => setQueueElement_start_req,
      start_ack => setQueueElement_start_ack,
      fin_req => setQueueElement_fin_req,
      fin_ack => setQueueElement_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(2 downto 2),
      accessMemory_call_acks => accessMemory_call_acks(2 downto 2),
      accessMemory_call_data => accessMemory_call_data(329 downto 220),
      accessMemory_call_tag => accessMemory_call_tag(5 downto 4),
      accessMemory_return_reqs => accessMemory_return_reqs(2 downto 2),
      accessMemory_return_acks => accessMemory_return_acks(2 downto 2),
      accessMemory_return_data => accessMemory_return_data(191 downto 128),
      accessMemory_return_tag => accessMemory_return_tag(5 downto 4),
      tag_in => setQueueElement_tag_in,
      tag_out => setQueueElement_tag_out-- 
    ); -- 
  -- module setQueuePointers
  setQueuePointers_q_base_address <= setQueuePointers_in_args(99 downto 64);
  setQueuePointers_wp <= setQueuePointers_in_args(63 downto 32);
  setQueuePointers_rp <= setQueuePointers_in_args(31 downto 0);
  -- call arbiter for module setQueuePointers
  setQueuePointers_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 2,
      call_data_width => 100,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => setQueuePointers_call_reqs,
      call_acks => setQueuePointers_call_acks,
      return_reqs => setQueuePointers_return_reqs,
      return_acks => setQueuePointers_return_acks,
      call_data  => setQueuePointers_call_data,
      call_tag  => setQueuePointers_call_tag,
      return_tag  => setQueuePointers_return_tag,
      call_mtag => setQueuePointers_tag_in,
      return_mtag => setQueuePointers_tag_out,
      call_mreq => setQueuePointers_start_req,
      call_mack => setQueuePointers_start_ack,
      return_mreq => setQueuePointers_fin_req,
      return_mack => setQueuePointers_fin_ack,
      call_mdata => setQueuePointers_in_args,
      clk => clk, 
      reset => reset --
    ); --
  setQueuePointers_instance:setQueuePointers-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => setQueuePointers_q_base_address,
      wp => setQueuePointers_wp,
      rp => setQueuePointers_rp,
      start_req => setQueuePointers_start_req,
      start_ack => setQueuePointers_start_ack,
      fin_req => setQueuePointers_fin_req,
      fin_ack => setQueuePointers_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(10 downto 10),
      accessMemory_call_acks => accessMemory_call_acks(10 downto 10),
      accessMemory_call_data => accessMemory_call_data(1209 downto 1100),
      accessMemory_call_tag => accessMemory_call_tag(21 downto 20),
      accessMemory_return_reqs => accessMemory_return_reqs(10 downto 10),
      accessMemory_return_acks => accessMemory_return_acks(10 downto 10),
      accessMemory_return_data => accessMemory_return_data(703 downto 640),
      accessMemory_return_tag => accessMemory_return_tag(21 downto 20),
      tag_in => setQueuePointers_tag_in,
      tag_out => setQueuePointers_tag_out-- 
    ); -- 
  -- module transmitEngineDaemon
  transmitEngineDaemon_instance:transmitEngineDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => transmitEngineDaemon_start_req,
      start_ack => transmitEngineDaemon_start_ack,
      fin_req => transmitEngineDaemon_fin_req,
      fin_ack => transmitEngineDaemon_fin_ack,
      clk => clk,
      reset => reset,
      FREE_Q => FREE_Q,
      LAST_READ_TX_QUEUE_INDEX => LAST_READ_TX_QUEUE_INDEX,
      CONTROL_REGISTER => CONTROL_REGISTER,
      NUMBER_OF_SERVERS => NUMBER_OF_SERVERS,
      LAST_READ_TX_QUEUE_INDEX_pipe_write_req => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(1 downto 0),
      LAST_READ_TX_QUEUE_INDEX_pipe_write_ack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(1 downto 0),
      LAST_READ_TX_QUEUE_INDEX_pipe_write_data => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(11 downto 0),
      AccessRegister_call_reqs => AccessRegister_call_reqs(0 downto 0),
      AccessRegister_call_acks => AccessRegister_call_acks(0 downto 0),
      AccessRegister_call_data => AccessRegister_call_data(42 downto 0),
      AccessRegister_call_tag => AccessRegister_call_tag(1 downto 0),
      AccessRegister_return_reqs => AccessRegister_return_reqs(0 downto 0),
      AccessRegister_return_acks => AccessRegister_return_acks(0 downto 0),
      AccessRegister_return_data => AccessRegister_return_data(31 downto 0),
      AccessRegister_return_tag => AccessRegister_return_tag(1 downto 0),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(0 downto 0),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(0 downto 0),
      pushIntoQueue_call_data => pushIntoQueue_call_data(68 downto 0),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(0 downto 0),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(0 downto 0),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(0 downto 0),
      pushIntoQueue_return_data => pushIntoQueue_return_data(0 downto 0),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(0 downto 0),
      getTxPacketPointerFromServer_call_reqs => getTxPacketPointerFromServer_call_reqs(0 downto 0),
      getTxPacketPointerFromServer_call_acks => getTxPacketPointerFromServer_call_acks(0 downto 0),
      getTxPacketPointerFromServer_call_data => getTxPacketPointerFromServer_call_data(5 downto 0),
      getTxPacketPointerFromServer_call_tag => getTxPacketPointerFromServer_call_tag(0 downto 0),
      getTxPacketPointerFromServer_return_reqs => getTxPacketPointerFromServer_return_reqs(0 downto 0),
      getTxPacketPointerFromServer_return_acks => getTxPacketPointerFromServer_return_acks(0 downto 0),
      getTxPacketPointerFromServer_return_data => getTxPacketPointerFromServer_return_data(32 downto 0),
      getTxPacketPointerFromServer_return_tag => getTxPacketPointerFromServer_return_tag(0 downto 0),
      transmitPacket_call_reqs => transmitPacket_call_reqs(0 downto 0),
      transmitPacket_call_acks => transmitPacket_call_acks(0 downto 0),
      transmitPacket_call_data => transmitPacket_call_data(31 downto 0),
      transmitPacket_call_tag => transmitPacket_call_tag(0 downto 0),
      transmitPacket_return_reqs => transmitPacket_return_reqs(0 downto 0),
      transmitPacket_return_acks => transmitPacket_return_acks(0 downto 0),
      transmitPacket_return_data => transmitPacket_return_data(0 downto 0),
      transmitPacket_return_tag => transmitPacket_return_tag(0 downto 0),
      tag_in => transmitEngineDaemon_tag_in,
      tag_out => transmitEngineDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  transmitEngineDaemon_tag_in <= (others => '0');
  transmitEngineDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => transmitEngineDaemon_start_req, start_ack => transmitEngineDaemon_start_ack,  fin_req => transmitEngineDaemon_fin_req,  fin_ack => transmitEngineDaemon_fin_ack);
  -- module transmitPacket
  transmitPacket_packet_pointer <= transmitPacket_in_args(31 downto 0);
  transmitPacket_out_args <= transmitPacket_status ;
  -- call arbiter for module transmitPacket
  transmitPacket_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 32,
      return_data_width => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => transmitPacket_call_reqs,
      call_acks => transmitPacket_call_acks,
      return_reqs => transmitPacket_return_reqs,
      return_acks => transmitPacket_return_acks,
      call_data  => transmitPacket_call_data,
      call_tag  => transmitPacket_call_tag,
      return_tag  => transmitPacket_return_tag,
      call_mtag => transmitPacket_tag_in,
      return_mtag => transmitPacket_tag_out,
      return_data =>transmitPacket_return_data,
      call_mreq => transmitPacket_start_req,
      call_mack => transmitPacket_start_ack,
      return_mreq => transmitPacket_fin_req,
      return_mack => transmitPacket_fin_ack,
      call_mdata => transmitPacket_in_args,
      return_mdata => transmitPacket_out_args,
      clk => clk, 
      reset => reset --
    ); --
  transmitPacket_instance:transmitPacket-- 
    generic map(tag_length => 2)
    port map(-- 
      packet_pointer => transmitPacket_packet_pointer,
      status => transmitPacket_status,
      start_req => transmitPacket_start_req,
      start_ack => transmitPacket_start_ack,
      fin_req => transmitPacket_fin_req,
      fin_ack => transmitPacket_fin_ack,
      clk => clk,
      reset => reset,
      nic_to_mac_transmit_pipe_pipe_write_req => nic_to_mac_transmit_pipe_pipe_write_req(1 downto 0),
      nic_to_mac_transmit_pipe_pipe_write_ack => nic_to_mac_transmit_pipe_pipe_write_ack(1 downto 0),
      nic_to_mac_transmit_pipe_pipe_write_data => nic_to_mac_transmit_pipe_pipe_write_data(145 downto 0),
      accessMemory_call_reqs => accessMemory_call_reqs(1 downto 0),
      accessMemory_call_acks => accessMemory_call_acks(1 downto 0),
      accessMemory_call_data => accessMemory_call_data(219 downto 0),
      accessMemory_call_tag => accessMemory_call_tag(3 downto 0),
      accessMemory_return_reqs => accessMemory_return_reqs(1 downto 0),
      accessMemory_return_acks => accessMemory_return_acks(1 downto 0),
      accessMemory_return_data => accessMemory_return_data(127 downto 0),
      accessMemory_return_tag => accessMemory_return_tag(3 downto 0),
      tag_in => transmitPacket_tag_in,
      tag_out => transmitPacket_tag_out-- 
    ); -- 
  -- module writeControlInformationToMem
  writeControlInformationToMem_base_buffer_pointer <= writeControlInformationToMem_in_args(51 downto 16);
  writeControlInformationToMem_packet_size <= writeControlInformationToMem_in_args(15 downto 8);
  writeControlInformationToMem_last_keep <= writeControlInformationToMem_in_args(7 downto 0);
  -- call arbiter for module writeControlInformationToMem
  writeControlInformationToMem_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 52,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeControlInformationToMem_call_reqs,
      call_acks => writeControlInformationToMem_call_acks,
      return_reqs => writeControlInformationToMem_return_reqs,
      return_acks => writeControlInformationToMem_return_acks,
      call_data  => writeControlInformationToMem_call_data,
      call_tag  => writeControlInformationToMem_call_tag,
      return_tag  => writeControlInformationToMem_return_tag,
      call_mtag => writeControlInformationToMem_tag_in,
      return_mtag => writeControlInformationToMem_tag_out,
      call_mreq => writeControlInformationToMem_start_req,
      call_mack => writeControlInformationToMem_start_ack,
      return_mreq => writeControlInformationToMem_fin_req,
      return_mack => writeControlInformationToMem_fin_ack,
      call_mdata => writeControlInformationToMem_in_args,
      clk => clk, 
      reset => reset --
    ); --
  writeControlInformationToMem_instance:writeControlInformationToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      base_buffer_pointer => writeControlInformationToMem_base_buffer_pointer,
      packet_size => writeControlInformationToMem_packet_size,
      last_keep => writeControlInformationToMem_last_keep,
      start_req => writeControlInformationToMem_start_req,
      start_ack => writeControlInformationToMem_start_ack,
      fin_req => writeControlInformationToMem_fin_req,
      fin_ack => writeControlInformationToMem_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(5 downto 5),
      accessMemory_call_acks => accessMemory_call_acks(5 downto 5),
      accessMemory_call_data => accessMemory_call_data(659 downto 550),
      accessMemory_call_tag => accessMemory_call_tag(11 downto 10),
      accessMemory_return_reqs => accessMemory_return_reqs(5 downto 5),
      accessMemory_return_acks => accessMemory_return_acks(5 downto 5),
      accessMemory_return_data => accessMemory_return_data(383 downto 320),
      accessMemory_return_tag => accessMemory_return_tag(11 downto 10),
      tag_in => writeControlInformationToMem_tag_in,
      tag_out => writeControlInformationToMem_tag_out-- 
    ); -- 
  -- module writeEthernetHeaderToMem
  writeEthernetHeaderToMem_buf_pointer <= writeEthernetHeaderToMem_in_args(35 downto 0);
  writeEthernetHeaderToMem_out_args <= writeEthernetHeaderToMem_buf_position ;
  -- call arbiter for module writeEthernetHeaderToMem
  writeEthernetHeaderToMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 36,
      return_data_width => 36,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeEthernetHeaderToMem_call_reqs,
      call_acks => writeEthernetHeaderToMem_call_acks,
      return_reqs => writeEthernetHeaderToMem_return_reqs,
      return_acks => writeEthernetHeaderToMem_return_acks,
      call_data  => writeEthernetHeaderToMem_call_data,
      call_tag  => writeEthernetHeaderToMem_call_tag,
      return_tag  => writeEthernetHeaderToMem_return_tag,
      call_mtag => writeEthernetHeaderToMem_tag_in,
      return_mtag => writeEthernetHeaderToMem_tag_out,
      return_data =>writeEthernetHeaderToMem_return_data,
      call_mreq => writeEthernetHeaderToMem_start_req,
      call_mack => writeEthernetHeaderToMem_start_ack,
      return_mreq => writeEthernetHeaderToMem_fin_req,
      return_mack => writeEthernetHeaderToMem_fin_ack,
      call_mdata => writeEthernetHeaderToMem_in_args,
      return_mdata => writeEthernetHeaderToMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  writeEthernetHeaderToMem_instance:writeEthernetHeaderToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      buf_pointer => writeEthernetHeaderToMem_buf_pointer,
      buf_position => writeEthernetHeaderToMem_buf_position,
      start_req => writeEthernetHeaderToMem_start_req,
      start_ack => writeEthernetHeaderToMem_start_ack,
      fin_req => writeEthernetHeaderToMem_fin_req,
      fin_ack => writeEthernetHeaderToMem_fin_ack,
      clk => clk,
      reset => reset,
      nic_rx_to_header_pipe_read_req => nic_rx_to_header_pipe_read_req(0 downto 0),
      nic_rx_to_header_pipe_read_ack => nic_rx_to_header_pipe_read_ack(0 downto 0),
      nic_rx_to_header_pipe_read_data => nic_rx_to_header_pipe_read_data(72 downto 0),
      accessMemory_call_reqs => accessMemory_call_reqs(4 downto 4),
      accessMemory_call_acks => accessMemory_call_acks(4 downto 4),
      accessMemory_call_data => accessMemory_call_data(549 downto 440),
      accessMemory_call_tag => accessMemory_call_tag(9 downto 8),
      accessMemory_return_reqs => accessMemory_return_reqs(4 downto 4),
      accessMemory_return_acks => accessMemory_return_acks(4 downto 4),
      accessMemory_return_data => accessMemory_return_data(319 downto 256),
      accessMemory_return_tag => accessMemory_return_tag(9 downto 8),
      tag_in => writeEthernetHeaderToMem_tag_in,
      tag_out => writeEthernetHeaderToMem_tag_out-- 
    ); -- 
  -- module writePayloadToMem
  writePayloadToMem_base_buf_pointer <= writePayloadToMem_in_args(71 downto 36);
  writePayloadToMem_buf_pointer <= writePayloadToMem_in_args(35 downto 0);
  writePayloadToMem_out_args <= writePayloadToMem_packet_size_32 & writePayloadToMem_bad_packet_identifier & writePayloadToMem_last_keep ;
  -- call arbiter for module writePayloadToMem
  writePayloadToMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 72,
      return_data_width => 17,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writePayloadToMem_call_reqs,
      call_acks => writePayloadToMem_call_acks,
      return_reqs => writePayloadToMem_return_reqs,
      return_acks => writePayloadToMem_return_acks,
      call_data  => writePayloadToMem_call_data,
      call_tag  => writePayloadToMem_call_tag,
      return_tag  => writePayloadToMem_return_tag,
      call_mtag => writePayloadToMem_tag_in,
      return_mtag => writePayloadToMem_tag_out,
      return_data =>writePayloadToMem_return_data,
      call_mreq => writePayloadToMem_start_req,
      call_mack => writePayloadToMem_start_ack,
      return_mreq => writePayloadToMem_fin_req,
      return_mack => writePayloadToMem_fin_ack,
      call_mdata => writePayloadToMem_in_args,
      return_mdata => writePayloadToMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  writePayloadToMem_instance:writePayloadToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      base_buf_pointer => writePayloadToMem_base_buf_pointer,
      buf_pointer => writePayloadToMem_buf_pointer,
      packet_size_32 => writePayloadToMem_packet_size_32,
      bad_packet_identifier => writePayloadToMem_bad_packet_identifier,
      last_keep => writePayloadToMem_last_keep,
      start_req => writePayloadToMem_start_req,
      start_ack => writePayloadToMem_start_ack,
      fin_req => writePayloadToMem_fin_req,
      fin_ack => writePayloadToMem_fin_ack,
      clk => clk,
      reset => reset,
      nic_rx_to_packet_pipe_read_req => nic_rx_to_packet_pipe_read_req(0 downto 0),
      nic_rx_to_packet_pipe_read_ack => nic_rx_to_packet_pipe_read_ack(0 downto 0),
      nic_rx_to_packet_pipe_read_data => nic_rx_to_packet_pipe_read_data(72 downto 0),
      accessMemory_call_reqs => accessMemory_call_reqs(3 downto 3),
      accessMemory_call_acks => accessMemory_call_acks(3 downto 3),
      accessMemory_call_data => accessMemory_call_data(439 downto 330),
      accessMemory_call_tag => accessMemory_call_tag(7 downto 6),
      accessMemory_return_reqs => accessMemory_return_reqs(3 downto 3),
      accessMemory_return_acks => accessMemory_return_acks(3 downto 3),
      accessMemory_return_data => accessMemory_return_data(255 downto 192),
      accessMemory_return_tag => accessMemory_return_tag(7 downto 6),
      tag_in => writePayloadToMem_tag_in,
      tag_out => writePayloadToMem_tag_out-- 
    ); -- 
  AFB_NIC_REQUEST_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe AFB_NIC_REQUEST",
      num_reads => 1,
      num_writes => 1,
      data_width => 74,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => AFB_NIC_REQUEST_pipe_read_req,
      read_ack => AFB_NIC_REQUEST_pipe_read_ack,
      read_data => AFB_NIC_REQUEST_pipe_read_data,
      write_req => AFB_NIC_REQUEST_pipe_write_req,
      write_ack => AFB_NIC_REQUEST_pipe_write_ack,
      write_data => AFB_NIC_REQUEST_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  AFB_NIC_RESPONSE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe AFB_NIC_RESPONSE",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => AFB_NIC_RESPONSE_pipe_read_req,
      read_ack => AFB_NIC_RESPONSE_pipe_read_ack,
      read_data => AFB_NIC_RESPONSE_pipe_read_data,
      write_req => AFB_NIC_RESPONSE_pipe_write_req,
      write_ack => AFB_NIC_RESPONSE_pipe_write_ack,
      write_data => AFB_NIC_RESPONSE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  CONTROL_REGISTER_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe CONTROL_REGISTER",
      volatile_flag => false,
      num_writes => 1,
      data_width => 32 --
    ) 
    port map( -- 
      read_data => CONTROL_REGISTER,
      write_req => CONTROL_REGISTER_pipe_write_req,
      write_ack => CONTROL_REGISTER_pipe_write_ack,
      write_data => CONTROL_REGISTER_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  FREE_Q_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe FREE_Q",
      volatile_flag => false,
      num_writes => 1,
      data_width => 36 --
    ) 
    port map( -- 
      read_data => FREE_Q,
      write_req => FREE_Q_pipe_write_req,
      write_ack => FREE_Q_pipe_write_ack,
      write_data => FREE_Q_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  LAST_READ_TX_QUEUE_INDEX_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe LAST_READ_TX_QUEUE_INDEX",
      volatile_flag => false,
      num_writes => 2,
      data_width => 6 --
    ) 
    port map( -- 
      read_data => LAST_READ_TX_QUEUE_INDEX,
      write_req => LAST_READ_TX_QUEUE_INDEX_pipe_write_req,
      write_ack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack,
      write_data => LAST_READ_TX_QUEUE_INDEX_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  LAST_WRITTEN_RX_QUEUE_INDEX_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe LAST_WRITTEN_RX_QUEUE_INDEX",
      volatile_flag => false,
      num_writes => 2,
      data_width => 6 --
    ) 
    port map( -- 
      read_data => LAST_WRITTEN_RX_QUEUE_INDEX,
      write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req,
      write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack,
      write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MEMORY_TO_NIC_RESPONSE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe MEMORY_TO_NIC_RESPONSE",
      num_reads => 1,
      num_writes => 1,
      data_width => 65,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => MEMORY_TO_NIC_RESPONSE_pipe_read_req,
      read_ack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack,
      read_data => MEMORY_TO_NIC_RESPONSE_pipe_read_data,
      write_req => MEMORY_TO_NIC_RESPONSE_pipe_write_req,
      write_ack => MEMORY_TO_NIC_RESPONSE_pipe_write_ack,
      write_data => MEMORY_TO_NIC_RESPONSE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_REQUEST_REGISTER_ACCESS_PIPE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_REQUEST_REGISTER_ACCESS_PIPE",
      num_reads => 1,
      num_writes => 1,
      data_width => 43,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req,
      read_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack,
      read_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data,
      write_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req,
      write_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack,
      write_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_RESPONSE_REGISTER_ACCESS_PIPE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_RESPONSE_REGISTER_ACCESS_PIPE",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req,
      read_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack,
      read_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data,
      write_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req,
      write_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack,
      write_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_TO_MEMORY_REQUEST_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_TO_MEMORY_REQUEST",
      num_reads => 1,
      num_writes => 1,
      data_width => 110,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => NIC_TO_MEMORY_REQUEST_pipe_read_req,
      read_ack => NIC_TO_MEMORY_REQUEST_pipe_read_ack,
      read_data => NIC_TO_MEMORY_REQUEST_pipe_read_data,
      write_req => NIC_TO_MEMORY_REQUEST_pipe_write_req,
      write_ack => NIC_TO_MEMORY_REQUEST_pipe_write_ack,
      write_data => NIC_TO_MEMORY_REQUEST_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NUMBER_OF_SERVERS_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe NUMBER_OF_SERVERS",
      volatile_flag => false,
      num_writes => 1,
      data_width => 32 --
    ) 
    port map( -- 
      read_data => NUMBER_OF_SERVERS,
      write_req => NUMBER_OF_SERVERS_pipe_write_req,
      write_ack => NUMBER_OF_SERVERS_pipe_write_ack,
      write_data => NUMBER_OF_SERVERS_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  mac_to_nic_data_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe mac_to_nic_data",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => mac_to_nic_data_pipe_read_req,
      read_ack => mac_to_nic_data_pipe_read_ack,
      read_data => mac_to_nic_data_pipe_read_data,
      write_req => mac_to_nic_data_pipe_write_req,
      write_ack => mac_to_nic_data_pipe_write_ack,
      write_data => mac_to_nic_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_rx_to_header_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_rx_to_header",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => nic_rx_to_header_pipe_read_req,
      read_ack => nic_rx_to_header_pipe_read_ack,
      read_data => nic_rx_to_header_pipe_read_data,
      write_req => nic_rx_to_header_pipe_write_req,
      write_ack => nic_rx_to_header_pipe_write_ack,
      write_data => nic_rx_to_header_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_rx_to_packet_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_rx_to_packet",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => nic_rx_to_packet_pipe_read_req,
      read_ack => nic_rx_to_packet_pipe_read_ack,
      read_data => nic_rx_to_packet_pipe_read_data,
      write_req => nic_rx_to_packet_pipe_write_req,
      write_ack => nic_rx_to_packet_pipe_write_ack,
      write_data => nic_rx_to_packet_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_to_mac_transmit_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_to_mac_transmit_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => nic_to_mac_transmit_pipe_pipe_read_req,
      read_ack => nic_to_mac_transmit_pipe_pipe_read_ack,
      read_data => nic_to_mac_transmit_pipe_pipe_read_data,
      write_req => nic_to_mac_transmit_pipe_pipe_write_req,
      write_ack => nic_to_mac_transmit_pipe_pipe_write_ack,
      write_data => nic_to_mac_transmit_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 2,
      num_stores => 1,
      addr_width => 6,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 6,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
